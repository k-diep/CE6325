* File: nand3.pex.sp
* Created: Fri Oct 27 14:55:11 2023
* Program "Calibre xRC"
* Version "v2013.2_18.13"
* 
.include "nand3.pex.sp.pex"
.subckt nand3  OUT VSS VDD A B C
* 
* C	C
* B	B
* A	A
* VDD	VDD
* VSS	VSS
* OUT	OUT
XD0_noxref N_VSS_D0_noxref_pos N_VDD_D0_noxref_neg DIODENWX  AREA=5.23258e-12
+ PERIM=9.15e-06
XMMN2 N_OUT_MMN2_d N_A_MMN2_g NET19 N_VSS_D0_noxref_pos NFET L=6.5e-08
+ W=5.6e-07 AD=1.8984e-13 AS=1.2796e-13 PD=1.798e-06 PS=1.017e-06 NRD=0.317857
+ NRS=0.408036 M=1 NF=1 CNR_SWITCH=1 PCCRIT=0 PAR=1 PTWELL=0 SA=3.39e-07
+ SB=1.158e-06 SD=0 PANW1=7.54e-15 PANW2=3.25e-15 PANW3=3.25e-15 PANW4=3.25e-15
+ PANW5=3.25e-15 PANW6=6.5e-15 PANW7=9.36e-15 PANW8=0 PANW9=0 PANW10=0
XMMN3 NET19 N_B_MMN3_g NET18 N_VSS_D0_noxref_pos NFET L=6.5e-08 W=5.6e-07
+ AD=1.2796e-13 AS=1.0192e-13 PD=1.017e-06 PS=9.24e-07 NRD=0.408036 NRS=0.325
+ M=1 NF=1 CNR_SWITCH=1 PCCRIT=0 PAR=1 PTWELL=0 SA=8.61e-07 SB=6.36e-07 SD=0
+ PANW1=7.54e-15 PANW2=3.25e-15 PANW3=3.25e-15 PANW4=3.25e-15 PANW5=3.25e-15
+ PANW6=6.5e-15 PANW7=9.36e-15 PANW8=0 PANW9=0 PANW10=0
XMMN0 NET18 N_C_MMN0_g N_VSS_MMN0_s N_VSS_D0_noxref_pos NFET L=6.5e-08
+ W=5.6e-07 AD=1.0192e-13 AS=1.1592e-13 PD=9.24e-07 PS=1.534e-06 NRD=0.325
+ NRS=0.178571 M=1 NF=1 CNR_SWITCH=1 PCCRIT=0 PAR=1 PTWELL=0 SA=1.29e-06
+ SB=2.07e-07 SD=0 PANW1=7.54e-15 PANW2=3.25e-15 PANW3=3.25e-15 PANW4=3.25e-15
+ PANW5=3.25e-15 PANW6=6.5e-15 PANW7=9.36e-15 PANW8=0 PANW9=0 PANW10=0
XMMP0 N_OUT_MMP0_d N_A_MMP0_g N_VDD_MMP0_s N_VDD_D0_noxref_neg PFET L=6.5e-08
+ W=9.6e-07 AD=2.1936e-13 AS=3.2544e-13 PD=1.417e-06 PS=2.598e-06 NRD=0.194792
+ NRS=0.185417 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=3.39e-07
+ SB=1.158e-06 SD=0 PANW1=0 PANW2=0 PANW3=1.885e-15 PANW4=3.25e-15
+ PANW5=3.25e-15 PANW6=6.5e-15 PANW7=7.54e-14 PANW8=1.5275e-14 PANW9=4.7515e-14
+ PANW10=9.6525e-14
XMMP3 N_OUT_MMP0_d N_B_MMP3_g N_VDD_MMP3_s N_VDD_D0_noxref_neg PFET L=6.5e-08
+ W=9.6e-07 AD=2.1936e-13 AS=1.7472e-13 PD=1.417e-06 PS=1.324e-06 NRD=0.28125
+ NRS=0.104167 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=8.61e-07
+ SB=6.36e-07 SD=0 PANW1=0 PANW2=0 PANW3=1.885e-15 PANW4=3.25e-15 PANW5=3.25e-15
+ PANW6=6.5e-15 PANW7=1.3e-14 PANW8=1.5275e-14 PANW9=1.72315e-13
+ PANW10=3.4125e-14
XMMP2 N_VDD_MMP3_s N_C_MMP2_g N_OUT_MMP2_s N_VDD_D0_noxref_neg PFET L=6.5e-08
+ W=9.6e-07 AD=1.7472e-13 AS=1.9872e-13 PD=1.324e-06 PS=2.334e-06 NRD=0.275
+ NRS=0.104167 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=1.29e-06
+ SB=2.07e-07 SD=0 PANW1=0 PANW2=0 PANW3=1.885e-15 PANW4=3.25e-15 PANW5=3.25e-15
+ PANW6=6.5e-15 PANW7=7.54e-14 PANW8=1.5275e-14 PANW9=4.7515e-14
+ PANW10=9.6525e-14
c_81 NET19 0 4.65971e-20
*
.include "nand3.pex.sp.NAND3.pxi"
*
.ends
*
*
