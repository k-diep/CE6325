module inv(in, out);
input in;
output out;
assign out = ~in;
endmodule

module nand2(a, b, out);
input a, b;
output out;
assign out = ~(a & b);
endmodule

module nand3(a, b, c, out);
input a, b, c;
output out;
assign out = ~(a & b & c);
endmodule

module nand4(a, b, c, d, out);
input a, b, c, d;
output out;
assign out = ~(a & b & c & d);
endmodule

module nor2(a, b, out);
input a, b;
output out;
assign out = ~(a | b);
endmodule

module nor3(a, b, c, out);
input a, b, c;
output out;
assign out = ~(a | b | c);
endmodule

module xor2(a, b, out);
input a, b;
output out;
assign out = (a ^ b);
endmodule

module aoi12(a, b, c, out);
input a, b, c;
output out;
assign out = ~(a | (b & c));
endmodule

module aoi22(a, b, c, d, out);
input a, b, c, d;
output out;
assign out = ~((a & b) | (c & d));
endmodule

module oai12(a, b, c, out);
input a, b, c;
output out;
assign out = ~(a & (b | c));
endmodule

module oai22(a, b, c, d, out);
input a, b, c, d;
output out;
assign out = ~((a | b) & (c | d));
endmodule

module dff( d, gclk, rnot, q);
input d, gclk, rnot;
output q;
reg q;
always @(posedge gclk or negedge rnot)
  if (rnot == 1'b0)
    q = 1'b0;
  else
    q = d;
endmodule


/////////////////////////////////////////////////////////////
// Created by: Synopsys DC Expert(TM) in wire load mode
// Version   : O-2018.06-SP1
// Date      : Sun Sep 24 14:31:30 2023
/////////////////////////////////////////////////////////////


module elevator ( requested_floor, destination_floor_elevator1, 
        destination_floor_elevator2, current_floor_elevator1, 
        current_floor_elevator2, clk, reset_elevator1, in_emergency_elevator1, 
        reset_elevator2, in_emergency_elevator2, direction_elevator1, 
        direction_elevator2, request_taken, elevator1_status, elevator2_status, 
        arrived_elevator1, arrived_elevator2, emergency_signal_elevator1, 
        emergency_signal_elevator2, current_floor_output_elevator1, 
        current_floor_output_elevator2, final_floor_elevator1, 
        final_floor_elevator2 );
  input [63:0] requested_floor;
  input [63:0] destination_floor_elevator1;
  input [63:0] destination_floor_elevator2;
  input [63:0] current_floor_elevator1;
  input [63:0] current_floor_elevator2;
  output [1:0] direction_elevator1;
  output [1:0] direction_elevator2;
  output [63:0] current_floor_output_elevator1;
  output [63:0] current_floor_output_elevator2;
  output [63:0] final_floor_elevator1;
  output [63:0] final_floor_elevator2;
  input clk, reset_elevator1, in_emergency_elevator1, reset_elevator2,
         in_emergency_elevator2;
  output request_taken, elevator1_status, elevator2_status, arrived_elevator1,
         arrived_elevator2, emergency_signal_elevator1,
         emergency_signal_elevator2;
  wire   N12, N13, N15, N16, N26, N27, N28, N29, N30, N31, N32, N33, N34, N35,
         N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46, N47, N48, N49,
         N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60, N61, N62, N63,
         N64, N65, N66, N67, N68, N69, N70, N71, N72, N73, N74, N75, N76, N77,
         N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88, N89, N90, N92,
         N93, N94, N95, N96, N97, N98, N99, N100, N101, N102, N103, N104, N105,
         N106, N107, N108, N109, N110, N111, N112, N113, N114, N115, N116,
         N117, N118, N119, N120, N121, N122, N123, N124, N125, N126, N127,
         N128, N129, N130, N131, N132, N133, N134, N135, N136, N137, N138,
         N139, N140, N141, N142, N143, N144, N145, N146, N147, N148, N149,
         N150, N151, N152, N153, N154, N156, N157, N158, N159, N160, N161,
         N162, N163, N164, N165, N166, N167, N168, N169, N170, N171, N172,
         N173, N174, N175, N176, N177, N178, N179, N180, N181, N182, N183,
         N184, N185, N186, N187, N188, N189, N190, N191, N192, N193, N194,
         N195, N196, N197, N198, N199, N200, N201, N202, N203, N204, N205,
         N206, N207, N208, N209, N210, N211, N212, N213, N214, N215, N216,
         N217, N218, N221, N223, N225, N230, N310, N311, N312, N313, N314,
         N315, N316, N317, N318, N319, N320, N321, N322, N323, N324, N325,
         N326, N327, N328, N329, N330, N331, N332, N333, N334, N335, N336,
         N337, N338, N339, N340, N341, N342, N343, N344, N345, N346, N347,
         N348, N349, N350, N351, N352, N353, N354, N355, N356, N357, N358,
         N359, N360, N361, N362, N363, N364, N365, N366, N367, N368, N369,
         N370, N371, N372, N373, N374, N376, N377, N378, N379, N380, N381,
         N382, N383, N384, N385, N386, N387, N388, N389, N390, N391, N392,
         N393, N394, N395, N396, N397, N398, N399, N400, N401, N402, N403,
         N404, N405, N406, N407, N408, N409, N410, N411, N412, N413, N414,
         N415, N416, N417, N418, N419, N420, N421, N422, N423, N424, N425,
         N426, N427, N428, N429, N430, N431, N432, N433, N434, N435, N436,
         N437, N438, N440, N441, N442, N443, N444, N445, N446, N447, N448,
         N449, N450, N451, N452, N453, N454, N455, N456, N457, N458, N459,
         N460, N461, N462, N463, N464, N465, N466, N467, N468, N469, N470,
         N471, N472, N473, N474, N475, N476, N477, N478, N479, N480, N481,
         N482, N483, N484, N485, N486, N487, N488, N489, N490, N491, N492,
         N493, N494, N495, N496, N497, N498, N499, N500, N501, N502, N505,
         N507, N509, N514, N604, N605, N606, N607, N609, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n32, n33, n34, n35, n36, n38,
         n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52,
         n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66,
         n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80,
         n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94,
         n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106,
         n107, n108, n109, n110, n111, n112, n113, n114, n115, n116, n117,
         n118, n119, n120, n121, n122, n123, n124, n125, n126, n127, n128,
         n129, n130, n131, n132, n133, n134, n135, n136, n137, n138, n139,
         n140, n141, n142, n143, n144, n145, n146, n147, n148, n149, n150,
         n151, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1165, n1166, n1167, n1168, n1169, n1170,
         n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180,
         n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190,
         n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200,
         n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210,
         n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220,
         n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230,
         n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240,
         n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250,
         n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260,
         n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270,
         n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280,
         n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290,
         n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300,
         n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310,
         n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320,
         n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330,
         n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340,
         n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350,
         n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360,
         n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370,
         n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380,
         n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390,
         n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400,
         n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410,
         n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420,
         n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430,
         \r126/SB , \r126/SA , \r125/SB , \r125/SA , \eq_47_3/SB ,
         \eq_47_3/SA , \eq_47_3/GT , \eq_47_3/LT , \ne_47/SB , \ne_47/SA ,
         \ne_47/EQ , \ne_47/GT , \ne_47/LT , \eq_42_3/SB , \eq_42_3/SA ,
         \eq_42_3/GT , \eq_42_3/LT , \ne_42/SA , \ne_42/EQ , \ne_42/GT ,
         \ne_42/LT , n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
         n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
         n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
         n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
         n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
         n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
         n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
         n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
         n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
         n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
         n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
         n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
         n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
         n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
         n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
         n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588,
         n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598,
         n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
         n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
         n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628,
         n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638,
         n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
         n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
         n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668,
         n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
         n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
         n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
         n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708,
         n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718,
         n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728,
         n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738,
         n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748,
         n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758,
         n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768,
         n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
         n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788,
         n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798,
         n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808,
         n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818,
         n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828,
         n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838,
         n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
         n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
         n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
         n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
         n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
         n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
         n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908,
         n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
         n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928,
         n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938,
         n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948,
         n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958,
         n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968,
         n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978,
         n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988,
         n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998,
         n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008,
         n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018,
         n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028,
         n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038,
         n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048,
         n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058,
         n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068,
         n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078,
         n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088,
         n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098,
         n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108,
         n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118,
         n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128,
         n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138,
         n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148,
         n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158,
         n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168,
         n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
         n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188,
         n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
         n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
         n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
         n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228,
         n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
         n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248,
         n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258,
         n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268,
         n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278,
         n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288,
         n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298,
         n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308,
         n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318,
         n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328,
         n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338,
         n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348,
         n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358,
         n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368,
         n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378,
         n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388,
         n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398,
         n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408,
         n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418,
         n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428,
         n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438,
         n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448,
         n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458,
         n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468,
         n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478,
         n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488,
         n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498,
         n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508,
         n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518,
         n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528,
         n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538,
         n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548,
         n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558,
         n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568,
         n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578,
         n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588,
         n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598,
         n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608,
         n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618,
         n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628,
         n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638,
         n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648,
         n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658,
         n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668,
         n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678,
         n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688,
         n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698,
         n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708,
         n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718,
         n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728,
         n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738,
         n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748,
         n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758,
         n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768,
         n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778,
         n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788,
         n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798,
         n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808,
         n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818,
         n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828,
         n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838,
         n2839, n2840, n2841, n2842;
  wire   [63:1] \r126/LTV2 ;
  wire   [63:1] \r126/LTV1 ;
  wire   [63:1] \r126/GTV2 ;
  wire   [63:1] \r126/GTV1 ;
  wire   [63:1] \r126/AEQB ;
  wire   [63:1] \r126/LTV ;
  wire   [63:1] \r126/GTV ;
  wire   [63:1] \r125/LTV2 ;
  wire   [63:1] \r125/LTV1 ;
  wire   [63:1] \r125/GTV2 ;
  wire   [63:1] \r125/GTV1 ;
  wire   [63:1] \r125/AEQB ;
  wire   [63:1] \r125/LTV ;
  wire   [63:1] \r125/GTV ;
  wire   [63:1] \eq_47_3/LTV2 ;
  wire   [63:1] \eq_47_3/LTV1 ;
  wire   [63:1] \eq_47_3/GTV2 ;
  wire   [63:1] \eq_47_3/GTV1 ;
  wire   [63:1] \eq_47_3/AEQB ;
  wire   [63:1] \eq_47_3/LTV ;
  wire   [63:1] \eq_47_3/GTV ;
  wire   [63:1] \ne_47/LTV2 ;
  wire   [63:1] \ne_47/LTV1 ;
  wire   [63:1] \ne_47/GTV2 ;
  wire   [63:1] \ne_47/GTV1 ;
  wire   [63:1] \ne_47/AEQB ;
  wire   [63:1] \ne_47/LTV ;
  wire   [63:1] \ne_47/GTV ;
  wire   [63:1] \eq_42_3/LTV2 ;
  wire   [63:1] \eq_42_3/LTV1 ;
  wire   [63:1] \eq_42_3/GTV2 ;
  wire   [63:1] \eq_42_3/GTV1 ;
  wire   [63:1] \eq_42_3/AEQB ;
  wire   [63:1] \eq_42_3/LTV ;
  wire   [63:1] \eq_42_3/GTV ;
  wire   [63:1] \ne_42/LTV2 ;
  wire   [63:1] \ne_42/LTV1 ;
  wire   [63:1] \ne_42/GTV2 ;
  wire   [63:1] \ne_42/GTV1 ;
  wire   [63:1] \ne_42/AEQB ;
  wire   [63:1] \ne_42/LTV ;
  wire   [63:1] \ne_42/GTV ;
  assign \eq_47_3/SB  = destination_floor_elevator2[63];
  assign current_floor_output_elevator2[63] = \eq_47_3/SA ;
  assign \ne_47/SB  = requested_floor[63];
  assign final_floor_elevator1[63] = \ne_47/SA ;
  assign \eq_42_3/SB  = destination_floor_elevator1[63];
  assign current_floor_output_elevator1[63] = \eq_42_3/SA ;
  assign final_floor_elevator2[63] = \ne_42/SA ;

  nand2 C2522 ( .a(n1511), .b(final_floor_elevator2[0]), .out(n1430) );
  nand2 C2521 ( .a(n1452), .b(N310), .out(n1429) );
  nand2 C2520 ( .a(n1429), .b(n1430), .out(N502) );
  nand2 C2518 ( .a(n1511), .b(final_floor_elevator2[1]), .out(n1428) );
  nand2 C2517 ( .a(n1451), .b(N311), .out(n1427) );
  nand2 C2516 ( .a(n1427), .b(n1428), .out(N501) );
  nand2 C2514 ( .a(n1511), .b(final_floor_elevator2[2]), .out(n1426) );
  nand2 C2513 ( .a(n1451), .b(N312), .out(n1425) );
  nand2 C2512 ( .a(n1425), .b(n1426), .out(N500) );
  nand2 C2510 ( .a(n1511), .b(final_floor_elevator2[3]), .out(n1424) );
  nand2 C2509 ( .a(n1451), .b(N313), .out(n1423) );
  nand2 C2508 ( .a(n1423), .b(n1424), .out(N499) );
  nand2 C2506 ( .a(n1511), .b(final_floor_elevator2[4]), .out(n1422) );
  nand2 C2505 ( .a(n1450), .b(N314), .out(n1421) );
  nand2 C2504 ( .a(n1421), .b(n1422), .out(N498) );
  nand2 C2502 ( .a(n1511), .b(final_floor_elevator2[5]), .out(n1420) );
  nand2 C2501 ( .a(n1450), .b(N315), .out(n1419) );
  nand2 C2500 ( .a(n1419), .b(n1420), .out(N497) );
  nand2 C2498 ( .a(n1510), .b(final_floor_elevator2[6]), .out(n1418) );
  nand2 C2497 ( .a(n1450), .b(N316), .out(n1417) );
  nand2 C2496 ( .a(n1417), .b(n1418), .out(N496) );
  nand2 C2494 ( .a(n1510), .b(final_floor_elevator2[7]), .out(n1416) );
  nand2 C2493 ( .a(n1449), .b(N317), .out(n1415) );
  nand2 C2492 ( .a(n1415), .b(n1416), .out(N495) );
  nand2 C2490 ( .a(n1510), .b(final_floor_elevator2[8]), .out(n1414) );
  nand2 C2489 ( .a(n1449), .b(N318), .out(n1413) );
  nand2 C2488 ( .a(n1413), .b(n1414), .out(N494) );
  nand2 C2486 ( .a(n1510), .b(final_floor_elevator2[9]), .out(n1412) );
  nand2 C2485 ( .a(n1449), .b(N319), .out(n1411) );
  nand2 C2484 ( .a(n1411), .b(n1412), .out(N493) );
  nand2 C2482 ( .a(n1510), .b(final_floor_elevator2[10]), .out(n1410) );
  nand2 C2481 ( .a(n1448), .b(N320), .out(n1409) );
  nand2 C2480 ( .a(n1409), .b(n1410), .out(N492) );
  nand2 C2478 ( .a(n1510), .b(final_floor_elevator2[11]), .out(n1408) );
  nand2 C2477 ( .a(n1448), .b(N321), .out(n1407) );
  nand2 C2476 ( .a(n1407), .b(n1408), .out(N491) );
  nand2 C2474 ( .a(n1510), .b(final_floor_elevator2[12]), .out(n1406) );
  nand2 C2473 ( .a(n1448), .b(N322), .out(n1405) );
  nand2 C2472 ( .a(n1405), .b(n1406), .out(N490) );
  nand2 C2470 ( .a(n1510), .b(final_floor_elevator2[13]), .out(n1404) );
  nand2 C2469 ( .a(n1447), .b(N323), .out(n1403) );
  nand2 C2468 ( .a(n1403), .b(n1404), .out(N489) );
  nand2 C2466 ( .a(n1510), .b(final_floor_elevator2[14]), .out(n1402) );
  nand2 C2465 ( .a(n1447), .b(N324), .out(n1401) );
  nand2 C2464 ( .a(n1401), .b(n1402), .out(N488) );
  nand2 C2462 ( .a(n1510), .b(final_floor_elevator2[15]), .out(n1400) );
  nand2 C2461 ( .a(n1447), .b(N325), .out(n1399) );
  nand2 C2460 ( .a(n1399), .b(n1400), .out(N487) );
  nand2 C2458 ( .a(n1510), .b(final_floor_elevator2[16]), .out(n1398) );
  nand2 C2457 ( .a(n1446), .b(N326), .out(n1397) );
  nand2 C2456 ( .a(n1397), .b(n1398), .out(N486) );
  nand2 C2454 ( .a(n1510), .b(final_floor_elevator2[17]), .out(n1396) );
  nand2 C2453 ( .a(n1446), .b(N327), .out(n1395) );
  nand2 C2452 ( .a(n1395), .b(n1396), .out(N485) );
  nand2 C2450 ( .a(n1509), .b(final_floor_elevator2[18]), .out(n1394) );
  nand2 C2449 ( .a(n1446), .b(N328), .out(n1393) );
  nand2 C2448 ( .a(n1393), .b(n1394), .out(N484) );
  nand2 C2446 ( .a(n1509), .b(final_floor_elevator2[19]), .out(n1392) );
  nand2 C2445 ( .a(n1445), .b(N329), .out(n1391) );
  nand2 C2444 ( .a(n1391), .b(n1392), .out(N483) );
  nand2 C2442 ( .a(n1509), .b(final_floor_elevator2[20]), .out(n1390) );
  nand2 C2441 ( .a(n1445), .b(N330), .out(n1389) );
  nand2 C2440 ( .a(n1389), .b(n1390), .out(N482) );
  nand2 C2438 ( .a(n1509), .b(final_floor_elevator2[21]), .out(n1388) );
  nand2 C2437 ( .a(n1445), .b(N331), .out(n1387) );
  nand2 C2436 ( .a(n1387), .b(n1388), .out(N481) );
  nand2 C2434 ( .a(n1509), .b(final_floor_elevator2[22]), .out(n1386) );
  nand2 C2433 ( .a(n1444), .b(N332), .out(n1385) );
  nand2 C2432 ( .a(n1385), .b(n1386), .out(N480) );
  nand2 C2430 ( .a(n1509), .b(final_floor_elevator2[23]), .out(n1384) );
  nand2 C2429 ( .a(n1444), .b(N333), .out(n1383) );
  nand2 C2428 ( .a(n1383), .b(n1384), .out(N479) );
  nand2 C2426 ( .a(n1509), .b(final_floor_elevator2[24]), .out(n1382) );
  nand2 C2425 ( .a(n1444), .b(N334), .out(n1381) );
  nand2 C2424 ( .a(n1381), .b(n1382), .out(N478) );
  nand2 C2422 ( .a(n1509), .b(final_floor_elevator2[25]), .out(n1380) );
  nand2 C2421 ( .a(n1443), .b(N335), .out(n1379) );
  nand2 C2420 ( .a(n1379), .b(n1380), .out(N477) );
  nand2 C2418 ( .a(n1509), .b(final_floor_elevator2[26]), .out(n1378) );
  nand2 C2417 ( .a(n1443), .b(N336), .out(n1377) );
  nand2 C2416 ( .a(n1377), .b(n1378), .out(N476) );
  nand2 C2414 ( .a(n1509), .b(final_floor_elevator2[27]), .out(n1376) );
  nand2 C2413 ( .a(n1443), .b(N337), .out(n1375) );
  nand2 C2412 ( .a(n1375), .b(n1376), .out(N475) );
  nand2 C2410 ( .a(n1509), .b(final_floor_elevator2[28]), .out(n1374) );
  nand2 C2409 ( .a(n1442), .b(N338), .out(n1373) );
  nand2 C2408 ( .a(n1373), .b(n1374), .out(N474) );
  nand2 C2406 ( .a(n1509), .b(final_floor_elevator2[29]), .out(n1372) );
  nand2 C2405 ( .a(n1442), .b(N339), .out(n1371) );
  nand2 C2404 ( .a(n1371), .b(n1372), .out(N473) );
  nand2 C2402 ( .a(n1508), .b(final_floor_elevator2[30]), .out(n1370) );
  nand2 C2401 ( .a(n1442), .b(N340), .out(n1369) );
  nand2 C2400 ( .a(n1369), .b(n1370), .out(N472) );
  nand2 C2398 ( .a(n1508), .b(final_floor_elevator2[31]), .out(n1368) );
  nand2 C2397 ( .a(n1441), .b(N341), .out(n1367) );
  nand2 C2396 ( .a(n1367), .b(n1368), .out(N471) );
  nand2 C2394 ( .a(n1508), .b(final_floor_elevator2[32]), .out(n1366) );
  nand2 C2393 ( .a(n1441), .b(N342), .out(n1365) );
  nand2 C2392 ( .a(n1365), .b(n1366), .out(N470) );
  nand2 C2390 ( .a(n1508), .b(final_floor_elevator2[33]), .out(n1364) );
  nand2 C2389 ( .a(n1441), .b(N343), .out(n1363) );
  nand2 C2388 ( .a(n1363), .b(n1364), .out(N469) );
  nand2 C2386 ( .a(n1508), .b(final_floor_elevator2[34]), .out(n1362) );
  nand2 C2385 ( .a(n1440), .b(N344), .out(n1361) );
  nand2 C2384 ( .a(n1361), .b(n1362), .out(N468) );
  nand2 C2382 ( .a(n1508), .b(final_floor_elevator2[35]), .out(n1360) );
  nand2 C2381 ( .a(n1440), .b(N345), .out(n1359) );
  nand2 C2380 ( .a(n1359), .b(n1360), .out(N467) );
  nand2 C2378 ( .a(n1508), .b(final_floor_elevator2[36]), .out(n1358) );
  nand2 C2377 ( .a(n1440), .b(N346), .out(n1357) );
  nand2 C2376 ( .a(n1357), .b(n1358), .out(N466) );
  nand2 C2374 ( .a(n1508), .b(final_floor_elevator2[37]), .out(n1356) );
  nand2 C2373 ( .a(n1439), .b(N347), .out(n1355) );
  nand2 C2372 ( .a(n1355), .b(n1356), .out(N465) );
  nand2 C2370 ( .a(n1508), .b(final_floor_elevator2[38]), .out(n1354) );
  nand2 C2369 ( .a(n1439), .b(N348), .out(n1353) );
  nand2 C2368 ( .a(n1353), .b(n1354), .out(N464) );
  nand2 C2366 ( .a(n1508), .b(final_floor_elevator2[39]), .out(n1352) );
  nand2 C2365 ( .a(n1439), .b(N349), .out(n1351) );
  nand2 C2364 ( .a(n1351), .b(n1352), .out(N463) );
  nand2 C2362 ( .a(n1508), .b(final_floor_elevator2[40]), .out(n1350) );
  nand2 C2361 ( .a(n1438), .b(N350), .out(n1349) );
  nand2 C2360 ( .a(n1349), .b(n1350), .out(N462) );
  nand2 C2358 ( .a(n1508), .b(final_floor_elevator2[41]), .out(n1348) );
  nand2 C2357 ( .a(n1438), .b(N351), .out(n1347) );
  nand2 C2356 ( .a(n1347), .b(n1348), .out(N461) );
  nand2 C2354 ( .a(n1507), .b(final_floor_elevator2[42]), .out(n1346) );
  nand2 C2353 ( .a(n1438), .b(N352), .out(n1345) );
  nand2 C2352 ( .a(n1345), .b(n1346), .out(N460) );
  nand2 C2350 ( .a(n1507), .b(final_floor_elevator2[43]), .out(n1344) );
  nand2 C2349 ( .a(n1437), .b(N353), .out(n1343) );
  nand2 C2348 ( .a(n1343), .b(n1344), .out(N459) );
  nand2 C2346 ( .a(n1507), .b(final_floor_elevator2[44]), .out(n1342) );
  nand2 C2345 ( .a(n1437), .b(N354), .out(n1341) );
  nand2 C2344 ( .a(n1341), .b(n1342), .out(N458) );
  nand2 C2342 ( .a(n1507), .b(final_floor_elevator2[45]), .out(n1340) );
  nand2 C2341 ( .a(n1437), .b(N355), .out(n1339) );
  nand2 C2340 ( .a(n1339), .b(n1340), .out(N457) );
  nand2 C2338 ( .a(n1507), .b(final_floor_elevator2[46]), .out(n1338) );
  nand2 C2337 ( .a(n1436), .b(N356), .out(n1337) );
  nand2 C2336 ( .a(n1337), .b(n1338), .out(N456) );
  nand2 C2334 ( .a(n1507), .b(final_floor_elevator2[47]), .out(n1336) );
  nand2 C2333 ( .a(n1436), .b(N357), .out(n1335) );
  nand2 C2332 ( .a(n1335), .b(n1336), .out(N455) );
  nand2 C2330 ( .a(n1507), .b(final_floor_elevator2[48]), .out(n1334) );
  nand2 C2329 ( .a(n1436), .b(N358), .out(n1333) );
  nand2 C2328 ( .a(n1333), .b(n1334), .out(N454) );
  nand2 C2326 ( .a(n1507), .b(final_floor_elevator2[49]), .out(n1332) );
  nand2 C2325 ( .a(n1435), .b(N359), .out(n1331) );
  nand2 C2324 ( .a(n1331), .b(n1332), .out(N453) );
  nand2 C2322 ( .a(n1512), .b(final_floor_elevator2[50]), .out(n1330) );
  nand2 C2321 ( .a(n1431), .b(N361), .out(n1329) );
  nand2 C2320 ( .a(n1329), .b(n1330), .out(N452) );
  nand2 C2318 ( .a(n1512), .b(final_floor_elevator2[51]), .out(n1328) );
  nand2 C2317 ( .a(n1431), .b(N362), .out(n1327) );
  nand2 C2316 ( .a(n1327), .b(n1328), .out(N451) );
  nand2 C2314 ( .a(n1512), .b(final_floor_elevator2[52]), .out(n1326) );
  nand2 C2313 ( .a(n1431), .b(N363), .out(n1325) );
  nand2 C2312 ( .a(n1325), .b(n1326), .out(N450) );
  nand2 C2310 ( .a(n1512), .b(final_floor_elevator2[53]), .out(n1324) );
  nand2 C2309 ( .a(n1432), .b(N364), .out(n1323) );
  nand2 C2308 ( .a(n1323), .b(n1324), .out(N449) );
  nand2 C2306 ( .a(n1512), .b(final_floor_elevator2[54]), .out(n1322) );
  nand2 C2305 ( .a(n1432), .b(N365), .out(n1321) );
  nand2 C2304 ( .a(n1321), .b(n1322), .out(N448) );
  nand2 C2302 ( .a(n1512), .b(final_floor_elevator2[55]), .out(n1320) );
  nand2 C2301 ( .a(n1432), .b(N366), .out(n1319) );
  nand2 C2300 ( .a(n1319), .b(n1320), .out(N447) );
  nand2 C2298 ( .a(n1512), .b(final_floor_elevator2[56]), .out(n1318) );
  nand2 C2297 ( .a(n1433), .b(N367), .out(n1317) );
  nand2 C2296 ( .a(n1317), .b(n1318), .out(N446) );
  nand2 C2294 ( .a(n1512), .b(final_floor_elevator2[57]), .out(n1316) );
  nand2 C2293 ( .a(n1433), .b(N368), .out(n1315) );
  nand2 C2292 ( .a(n1315), .b(n1316), .out(N445) );
  nand2 C2290 ( .a(n1511), .b(final_floor_elevator2[58]), .out(n1314) );
  nand2 C2289 ( .a(n1433), .b(N369), .out(n1313) );
  nand2 C2288 ( .a(n1313), .b(n1314), .out(N444) );
  nand2 C2286 ( .a(n1511), .b(final_floor_elevator2[59]), .out(n1312) );
  nand2 C2285 ( .a(n1434), .b(N370), .out(n1311) );
  nand2 C2284 ( .a(n1311), .b(n1312), .out(N443) );
  nand2 C2282 ( .a(n1511), .b(final_floor_elevator2[60]), .out(n1310) );
  nand2 C2281 ( .a(n1434), .b(N371), .out(n1309) );
  nand2 C2280 ( .a(n1309), .b(n1310), .out(N442) );
  nand2 C2278 ( .a(n1511), .b(final_floor_elevator2[61]), .out(n1308) );
  nand2 C2277 ( .a(n1434), .b(N372), .out(n1307) );
  nand2 C2276 ( .a(n1307), .b(n1308), .out(N441) );
  nand2 C2274 ( .a(n1511), .b(final_floor_elevator2[62]), .out(n1306) );
  nand2 C2273 ( .a(n1435), .b(N373), .out(n1305) );
  nand2 C2272 ( .a(n1305), .b(n1306), .out(N440) );
  nand2 C2270 ( .a(n1511), .b(\ne_42/SA ), .out(n1304) );
  nand2 C2269 ( .a(n1435), .b(N374), .out(n1303) );
  nand2 C2268 ( .a(n1303), .b(n1304), .out(\r126/SA ) );
  nand2 C2266 ( .a(n1639), .b(current_floor_output_elevator2[0]), .out(n647)
         );
  nand2 C2265 ( .a(n1611), .b(current_floor_elevator2[0]), .out(n646) );
  nand2 C2262 ( .a(n1639), .b(current_floor_output_elevator2[1]), .out(n643)
         );
  nand2 C2261 ( .a(n1611), .b(current_floor_elevator2[1]), .out(n642) );
  nand2 C2258 ( .a(n1639), .b(current_floor_output_elevator2[2]), .out(n645)
         );
  nand2 C2257 ( .a(n1611), .b(current_floor_elevator2[2]), .out(n644) );
  nand2 C2254 ( .a(n1638), .b(current_floor_output_elevator2[3]), .out(n649)
         );
  nand2 C2253 ( .a(n1610), .b(current_floor_elevator2[3]), .out(n648) );
  nand2 C2250 ( .a(n1638), .b(current_floor_output_elevator2[4]), .out(n651)
         );
  nand2 C2249 ( .a(n1610), .b(current_floor_elevator2[4]), .out(n650) );
  nand2 C2246 ( .a(n1638), .b(current_floor_output_elevator2[5]), .out(n653)
         );
  nand2 C2245 ( .a(n1610), .b(current_floor_elevator2[5]), .out(n652) );
  nand2 C2242 ( .a(n1637), .b(current_floor_output_elevator2[6]), .out(n655)
         );
  nand2 C2241 ( .a(n1610), .b(current_floor_elevator2[6]), .out(n654) );
  nand2 C2238 ( .a(n1637), .b(current_floor_output_elevator2[7]), .out(n657)
         );
  nand2 C2237 ( .a(n1610), .b(current_floor_elevator2[7]), .out(n656) );
  nand2 C2234 ( .a(n1637), .b(current_floor_output_elevator2[8]), .out(n659)
         );
  nand2 C2233 ( .a(n1610), .b(current_floor_elevator2[8]), .out(n658) );
  nand2 C2230 ( .a(n1636), .b(current_floor_output_elevator2[9]), .out(n661)
         );
  nand2 C2229 ( .a(n1610), .b(current_floor_elevator2[9]), .out(n660) );
  nand2 C2226 ( .a(n1636), .b(current_floor_output_elevator2[10]), .out(n663)
         );
  nand2 C2225 ( .a(n1610), .b(current_floor_elevator2[10]), .out(n662) );
  nand2 C2222 ( .a(n1636), .b(current_floor_output_elevator2[11]), .out(n665)
         );
  nand2 C2221 ( .a(n1610), .b(current_floor_elevator2[11]), .out(n664) );
  nand2 C2218 ( .a(n1635), .b(current_floor_output_elevator2[12]), .out(n667)
         );
  nand2 C2217 ( .a(n1610), .b(current_floor_elevator2[12]), .out(n666) );
  nand2 C2214 ( .a(n1635), .b(current_floor_output_elevator2[13]), .out(n669)
         );
  nand2 C2213 ( .a(n1610), .b(current_floor_elevator2[13]), .out(n668) );
  nand2 C2210 ( .a(n1635), .b(current_floor_output_elevator2[14]), .out(n671)
         );
  nand2 C2209 ( .a(n1610), .b(current_floor_elevator2[14]), .out(n670) );
  nand2 C2206 ( .a(n1634), .b(current_floor_output_elevator2[15]), .out(n673)
         );
  nand2 C2205 ( .a(n1609), .b(current_floor_elevator2[15]), .out(n672) );
  nand2 C2202 ( .a(n1634), .b(current_floor_output_elevator2[16]), .out(n675)
         );
  nand2 C2201 ( .a(n1609), .b(current_floor_elevator2[16]), .out(n674) );
  nand2 C2198 ( .a(n1634), .b(current_floor_output_elevator2[17]), .out(n677)
         );
  nand2 C2197 ( .a(n1609), .b(current_floor_elevator2[17]), .out(n676) );
  nand2 C2194 ( .a(n1633), .b(current_floor_output_elevator2[18]), .out(n679)
         );
  nand2 C2193 ( .a(n1609), .b(current_floor_elevator2[18]), .out(n678) );
  nand2 C2190 ( .a(n1633), .b(current_floor_output_elevator2[19]), .out(n681)
         );
  nand2 C2189 ( .a(n1609), .b(current_floor_elevator2[19]), .out(n680) );
  nand2 C2186 ( .a(n1633), .b(current_floor_output_elevator2[20]), .out(n683)
         );
  nand2 C2185 ( .a(n1609), .b(current_floor_elevator2[20]), .out(n682) );
  nand2 C2182 ( .a(n1632), .b(current_floor_output_elevator2[21]), .out(n685)
         );
  nand2 C2181 ( .a(n1609), .b(current_floor_elevator2[21]), .out(n684) );
  nand2 C2178 ( .a(n1632), .b(current_floor_output_elevator2[22]), .out(n687)
         );
  nand2 C2177 ( .a(n1609), .b(current_floor_elevator2[22]), .out(n686) );
  nand2 C2174 ( .a(n1632), .b(current_floor_output_elevator2[23]), .out(n689)
         );
  nand2 C2173 ( .a(n1609), .b(current_floor_elevator2[23]), .out(n688) );
  nand2 C2170 ( .a(n1631), .b(current_floor_output_elevator2[24]), .out(n691)
         );
  nand2 C2169 ( .a(n1609), .b(current_floor_elevator2[24]), .out(n690) );
  nand2 C2166 ( .a(n1631), .b(current_floor_output_elevator2[25]), .out(n693)
         );
  nand2 C2165 ( .a(n1609), .b(current_floor_elevator2[25]), .out(n692) );
  nand2 C2162 ( .a(n1631), .b(current_floor_output_elevator2[26]), .out(n695)
         );
  nand2 C2161 ( .a(n1609), .b(current_floor_elevator2[26]), .out(n694) );
  nand2 C2158 ( .a(n1630), .b(current_floor_output_elevator2[27]), .out(n697)
         );
  nand2 C2157 ( .a(n1608), .b(current_floor_elevator2[27]), .out(n696) );
  nand2 C2154 ( .a(n1630), .b(current_floor_output_elevator2[28]), .out(n699)
         );
  nand2 C2153 ( .a(n1608), .b(current_floor_elevator2[28]), .out(n698) );
  nand2 C2150 ( .a(n1630), .b(current_floor_output_elevator2[29]), .out(n701)
         );
  nand2 C2149 ( .a(n1608), .b(current_floor_elevator2[29]), .out(n700) );
  nand2 C2146 ( .a(n1629), .b(current_floor_output_elevator2[30]), .out(n703)
         );
  nand2 C2145 ( .a(n1608), .b(current_floor_elevator2[30]), .out(n702) );
  nand2 C2142 ( .a(n1629), .b(current_floor_output_elevator2[31]), .out(n705)
         );
  nand2 C2141 ( .a(n1608), .b(current_floor_elevator2[31]), .out(n704) );
  nand2 C2138 ( .a(n1629), .b(current_floor_output_elevator2[32]), .out(n707)
         );
  nand2 C2137 ( .a(n1608), .b(current_floor_elevator2[32]), .out(n706) );
  nand2 C2134 ( .a(n1628), .b(current_floor_output_elevator2[33]), .out(n709)
         );
  nand2 C2133 ( .a(n1608), .b(current_floor_elevator2[33]), .out(n708) );
  nand2 C2130 ( .a(n1628), .b(current_floor_output_elevator2[34]), .out(n711)
         );
  nand2 C2129 ( .a(n1608), .b(current_floor_elevator2[34]), .out(n710) );
  nand2 C2126 ( .a(n1628), .b(current_floor_output_elevator2[35]), .out(n713)
         );
  nand2 C2125 ( .a(n1608), .b(current_floor_elevator2[35]), .out(n712) );
  nand2 C2122 ( .a(n1627), .b(current_floor_output_elevator2[36]), .out(n715)
         );
  nand2 C2121 ( .a(n1608), .b(current_floor_elevator2[36]), .out(n714) );
  nand2 C2118 ( .a(n1627), .b(current_floor_output_elevator2[37]), .out(n717)
         );
  nand2 C2117 ( .a(n1608), .b(current_floor_elevator2[37]), .out(n716) );
  nand2 C2114 ( .a(n1627), .b(current_floor_output_elevator2[38]), .out(n719)
         );
  nand2 C2113 ( .a(n1608), .b(current_floor_elevator2[38]), .out(n718) );
  nand2 C2110 ( .a(n1626), .b(current_floor_output_elevator2[39]), .out(n721)
         );
  nand2 C2109 ( .a(n1607), .b(current_floor_elevator2[39]), .out(n720) );
  nand2 C2106 ( .a(n1626), .b(current_floor_output_elevator2[40]), .out(n723)
         );
  nand2 C2105 ( .a(n1607), .b(current_floor_elevator2[40]), .out(n722) );
  nand2 C2102 ( .a(n1626), .b(current_floor_output_elevator2[41]), .out(n725)
         );
  nand2 C2101 ( .a(n1607), .b(current_floor_elevator2[41]), .out(n724) );
  nand2 C2098 ( .a(n1625), .b(current_floor_output_elevator2[42]), .out(n727)
         );
  nand2 C2097 ( .a(n1607), .b(current_floor_elevator2[42]), .out(n726) );
  nand2 C2094 ( .a(n1625), .b(current_floor_output_elevator2[43]), .out(n729)
         );
  nand2 C2093 ( .a(n1607), .b(current_floor_elevator2[43]), .out(n728) );
  nand2 C2090 ( .a(n1625), .b(current_floor_output_elevator2[44]), .out(n731)
         );
  nand2 C2089 ( .a(n1607), .b(current_floor_elevator2[44]), .out(n730) );
  nand2 C2086 ( .a(n1624), .b(current_floor_output_elevator2[45]), .out(n733)
         );
  nand2 C2085 ( .a(n1607), .b(current_floor_elevator2[45]), .out(n732) );
  nand2 C2082 ( .a(n1624), .b(current_floor_output_elevator2[46]), .out(n735)
         );
  nand2 C2081 ( .a(n1607), .b(current_floor_elevator2[46]), .out(n734) );
  nand2 C2078 ( .a(n1624), .b(current_floor_output_elevator2[47]), .out(n737)
         );
  nand2 C2077 ( .a(n1607), .b(current_floor_elevator2[47]), .out(n736) );
  nand2 C2074 ( .a(n1623), .b(current_floor_output_elevator2[48]), .out(n739)
         );
  nand2 C2073 ( .a(n1607), .b(current_floor_elevator2[48]), .out(n738) );
  nand2 C2070 ( .a(n1623), .b(current_floor_output_elevator2[49]), .out(n741)
         );
  nand2 C2069 ( .a(n1607), .b(current_floor_elevator2[49]), .out(n740) );
  nand2 C2066 ( .a(n1623), .b(current_floor_output_elevator2[50]), .out(n743)
         );
  nand2 C2065 ( .a(n1607), .b(current_floor_elevator2[50]), .out(n742) );
  nand2 C2062 ( .a(n1622), .b(current_floor_output_elevator2[51]), .out(n745)
         );
  nand2 C2061 ( .a(n1606), .b(current_floor_elevator2[51]), .out(n744) );
  nand2 C2058 ( .a(n1622), .b(current_floor_output_elevator2[52]), .out(n747)
         );
  nand2 C2057 ( .a(n1606), .b(current_floor_elevator2[52]), .out(n746) );
  nand2 C2054 ( .a(n1622), .b(current_floor_output_elevator2[53]), .out(n749)
         );
  nand2 C2053 ( .a(n1606), .b(current_floor_elevator2[53]), .out(n748) );
  nand2 C2050 ( .a(n1621), .b(current_floor_output_elevator2[54]), .out(n751)
         );
  nand2 C2049 ( .a(n1606), .b(current_floor_elevator2[54]), .out(n750) );
  nand2 C2046 ( .a(n1621), .b(current_floor_output_elevator2[55]), .out(n753)
         );
  nand2 C2045 ( .a(n1606), .b(current_floor_elevator2[55]), .out(n752) );
  nand2 C2042 ( .a(n1621), .b(current_floor_output_elevator2[56]), .out(n755)
         );
  nand2 C2041 ( .a(n1606), .b(current_floor_elevator2[56]), .out(n754) );
  nand2 C2038 ( .a(n1620), .b(current_floor_output_elevator2[57]), .out(n757)
         );
  nand2 C2037 ( .a(n1606), .b(current_floor_elevator2[57]), .out(n756) );
  nand2 C2034 ( .a(n1620), .b(current_floor_output_elevator2[58]), .out(n759)
         );
  nand2 C2033 ( .a(n1606), .b(current_floor_elevator2[58]), .out(n758) );
  nand2 C2030 ( .a(n1620), .b(current_floor_output_elevator2[59]), .out(n761)
         );
  nand2 C2029 ( .a(n1606), .b(current_floor_elevator2[59]), .out(n760) );
  nand2 C2026 ( .a(n1619), .b(current_floor_output_elevator2[60]), .out(n763)
         );
  nand2 C2025 ( .a(n1606), .b(current_floor_elevator2[60]), .out(n762) );
  nand2 C2022 ( .a(n1619), .b(current_floor_output_elevator2[61]), .out(n765)
         );
  nand2 C2021 ( .a(n1606), .b(current_floor_elevator2[61]), .out(n764) );
  nand2 C2018 ( .a(n1619), .b(current_floor_output_elevator2[62]), .out(n767)
         );
  nand2 C2017 ( .a(n1606), .b(current_floor_elevator2[62]), .out(n766) );
  nand2 C2014 ( .a(n1618), .b(\eq_47_3/SA ), .out(n769) );
  nand2 C2013 ( .a(n1605), .b(current_floor_elevator2[63]), .out(n768) );
  nand2 C1996 ( .a(n1593), .b(final_floor_elevator1[0]), .out(n1302) );
  nand2 C1995 ( .a(n1534), .b(N26), .out(n1301) );
  nand2 C1994 ( .a(n1301), .b(n1302), .out(N218) );
  nand2 C1992 ( .a(n1593), .b(final_floor_elevator1[1]), .out(n1300) );
  nand2 C1991 ( .a(n1533), .b(N27), .out(n1299) );
  nand2 C1990 ( .a(n1299), .b(n1300), .out(N217) );
  nand2 C1988 ( .a(n1593), .b(final_floor_elevator1[2]), .out(n1298) );
  nand2 C1987 ( .a(n1533), .b(N28), .out(n1297) );
  nand2 C1986 ( .a(n1297), .b(n1298), .out(N216) );
  nand2 C1984 ( .a(n1593), .b(final_floor_elevator1[3]), .out(n1296) );
  nand2 C1983 ( .a(n1533), .b(N29), .out(n1295) );
  nand2 C1982 ( .a(n1295), .b(n1296), .out(N215) );
  nand2 C1980 ( .a(n1593), .b(final_floor_elevator1[4]), .out(n1294) );
  nand2 C1979 ( .a(n1532), .b(N30), .out(n1293) );
  nand2 C1978 ( .a(n1293), .b(n1294), .out(N214) );
  nand2 C1976 ( .a(n1593), .b(final_floor_elevator1[5]), .out(n1292) );
  nand2 C1975 ( .a(n1532), .b(N31), .out(n1291) );
  nand2 C1974 ( .a(n1291), .b(n1292), .out(N213) );
  nand2 C1972 ( .a(n1593), .b(final_floor_elevator1[6]), .out(n1290) );
  nand2 C1971 ( .a(n1532), .b(N32), .out(n1289) );
  nand2 C1970 ( .a(n1289), .b(n1290), .out(N212) );
  nand2 C1968 ( .a(n1592), .b(final_floor_elevator1[7]), .out(n1288) );
  nand2 C1967 ( .a(n1531), .b(N33), .out(n1287) );
  nand2 C1966 ( .a(n1287), .b(n1288), .out(N211) );
  nand2 C1964 ( .a(n1592), .b(final_floor_elevator1[8]), .out(n1286) );
  nand2 C1963 ( .a(n1531), .b(N34), .out(n1285) );
  nand2 C1962 ( .a(n1285), .b(n1286), .out(N210) );
  nand2 C1960 ( .a(n1592), .b(final_floor_elevator1[9]), .out(n1284) );
  nand2 C1959 ( .a(n1531), .b(N35), .out(n1283) );
  nand2 C1958 ( .a(n1283), .b(n1284), .out(N209) );
  nand2 C1956 ( .a(n1592), .b(final_floor_elevator1[10]), .out(n1282) );
  nand2 C1955 ( .a(n1530), .b(N36), .out(n1281) );
  nand2 C1954 ( .a(n1281), .b(n1282), .out(N208) );
  nand2 C1952 ( .a(n1592), .b(final_floor_elevator1[11]), .out(n1280) );
  nand2 C1951 ( .a(n1530), .b(N37), .out(n1279) );
  nand2 C1950 ( .a(n1279), .b(n1280), .out(N207) );
  nand2 C1948 ( .a(n1592), .b(final_floor_elevator1[12]), .out(n1278) );
  nand2 C1947 ( .a(n1530), .b(N38), .out(n1277) );
  nand2 C1946 ( .a(n1277), .b(n1278), .out(N206) );
  nand2 C1944 ( .a(n1592), .b(final_floor_elevator1[13]), .out(n1276) );
  nand2 C1943 ( .a(n1529), .b(N39), .out(n1275) );
  nand2 C1942 ( .a(n1275), .b(n1276), .out(N205) );
  nand2 C1940 ( .a(n1592), .b(final_floor_elevator1[14]), .out(n1274) );
  nand2 C1939 ( .a(n1529), .b(N40), .out(n1273) );
  nand2 C1938 ( .a(n1273), .b(n1274), .out(N204) );
  nand2 C1936 ( .a(n1592), .b(final_floor_elevator1[15]), .out(n1272) );
  nand2 C1935 ( .a(n1529), .b(N41), .out(n1271) );
  nand2 C1934 ( .a(n1271), .b(n1272), .out(N203) );
  nand2 C1932 ( .a(n1592), .b(final_floor_elevator1[16]), .out(n1270) );
  nand2 C1931 ( .a(n1528), .b(N42), .out(n1269) );
  nand2 C1930 ( .a(n1269), .b(n1270), .out(N202) );
  nand2 C1928 ( .a(n1592), .b(final_floor_elevator1[17]), .out(n1268) );
  nand2 C1927 ( .a(n1528), .b(N43), .out(n1267) );
  nand2 C1926 ( .a(n1267), .b(n1268), .out(N201) );
  nand2 C1924 ( .a(n1592), .b(final_floor_elevator1[18]), .out(n1266) );
  nand2 C1923 ( .a(n1528), .b(N44), .out(n1265) );
  nand2 C1922 ( .a(n1265), .b(n1266), .out(N200) );
  nand2 C1920 ( .a(n1591), .b(final_floor_elevator1[19]), .out(n1264) );
  nand2 C1919 ( .a(n1527), .b(N45), .out(n1263) );
  nand2 C1918 ( .a(n1263), .b(n1264), .out(N199) );
  nand2 C1916 ( .a(n1591), .b(final_floor_elevator1[20]), .out(n1262) );
  nand2 C1915 ( .a(n1527), .b(N46), .out(n1261) );
  nand2 C1914 ( .a(n1261), .b(n1262), .out(N198) );
  nand2 C1912 ( .a(n1591), .b(final_floor_elevator1[21]), .out(n1260) );
  nand2 C1911 ( .a(n1527), .b(N47), .out(n1259) );
  nand2 C1910 ( .a(n1259), .b(n1260), .out(N197) );
  nand2 C1908 ( .a(n1591), .b(final_floor_elevator1[22]), .out(n1258) );
  nand2 C1907 ( .a(n1526), .b(N48), .out(n1257) );
  nand2 C1906 ( .a(n1257), .b(n1258), .out(N196) );
  nand2 C1904 ( .a(n1591), .b(final_floor_elevator1[23]), .out(n1256) );
  nand2 C1903 ( .a(n1526), .b(N49), .out(n1255) );
  nand2 C1902 ( .a(n1255), .b(n1256), .out(N195) );
  nand2 C1900 ( .a(n1591), .b(final_floor_elevator1[24]), .out(n1254) );
  nand2 C1899 ( .a(n1526), .b(N50), .out(n1253) );
  nand2 C1898 ( .a(n1253), .b(n1254), .out(N194) );
  nand2 C1896 ( .a(n1591), .b(final_floor_elevator1[25]), .out(n1252) );
  nand2 C1895 ( .a(n1525), .b(N51), .out(n1251) );
  nand2 C1894 ( .a(n1251), .b(n1252), .out(N193) );
  nand2 C1892 ( .a(n1591), .b(final_floor_elevator1[26]), .out(n1250) );
  nand2 C1891 ( .a(n1525), .b(N52), .out(n1249) );
  nand2 C1890 ( .a(n1249), .b(n1250), .out(N192) );
  nand2 C1888 ( .a(n1591), .b(final_floor_elevator1[27]), .out(n1248) );
  nand2 C1887 ( .a(n1525), .b(N53), .out(n1247) );
  nand2 C1886 ( .a(n1247), .b(n1248), .out(N191) );
  nand2 C1884 ( .a(n1591), .b(final_floor_elevator1[28]), .out(n1246) );
  nand2 C1883 ( .a(n1524), .b(N54), .out(n1245) );
  nand2 C1882 ( .a(n1245), .b(n1246), .out(N190) );
  nand2 C1880 ( .a(n1591), .b(final_floor_elevator1[29]), .out(n1244) );
  nand2 C1879 ( .a(n1524), .b(N55), .out(n1243) );
  nand2 C1878 ( .a(n1243), .b(n1244), .out(N189) );
  nand2 C1876 ( .a(n1591), .b(final_floor_elevator1[30]), .out(n1242) );
  nand2 C1875 ( .a(n1524), .b(N56), .out(n1241) );
  nand2 C1874 ( .a(n1241), .b(n1242), .out(N188) );
  nand2 C1872 ( .a(n1590), .b(final_floor_elevator1[31]), .out(n1240) );
  nand2 C1871 ( .a(n1523), .b(N57), .out(n1239) );
  nand2 C1870 ( .a(n1239), .b(n1240), .out(N187) );
  nand2 C1868 ( .a(n1590), .b(final_floor_elevator1[32]), .out(n1238) );
  nand2 C1867 ( .a(n1523), .b(N58), .out(n1237) );
  nand2 C1866 ( .a(n1237), .b(n1238), .out(N186) );
  nand2 C1864 ( .a(n1590), .b(final_floor_elevator1[33]), .out(n1236) );
  nand2 C1863 ( .a(n1523), .b(N59), .out(n1235) );
  nand2 C1862 ( .a(n1235), .b(n1236), .out(N185) );
  nand2 C1860 ( .a(n1590), .b(final_floor_elevator1[34]), .out(n1234) );
  nand2 C1859 ( .a(n1522), .b(N60), .out(n1233) );
  nand2 C1858 ( .a(n1233), .b(n1234), .out(N184) );
  nand2 C1856 ( .a(n1590), .b(final_floor_elevator1[35]), .out(n1232) );
  nand2 C1855 ( .a(n1522), .b(N61), .out(n1231) );
  nand2 C1854 ( .a(n1231), .b(n1232), .out(N183) );
  nand2 C1852 ( .a(n1590), .b(final_floor_elevator1[36]), .out(n1230) );
  nand2 C1851 ( .a(n1522), .b(N62), .out(n1229) );
  nand2 C1850 ( .a(n1229), .b(n1230), .out(N182) );
  nand2 C1848 ( .a(n1590), .b(final_floor_elevator1[37]), .out(n1228) );
  nand2 C1847 ( .a(n1521), .b(N63), .out(n1227) );
  nand2 C1846 ( .a(n1227), .b(n1228), .out(N181) );
  nand2 C1844 ( .a(n1590), .b(final_floor_elevator1[38]), .out(n1226) );
  nand2 C1843 ( .a(n1521), .b(N64), .out(n1225) );
  nand2 C1842 ( .a(n1225), .b(n1226), .out(N180) );
  nand2 C1840 ( .a(n1590), .b(final_floor_elevator1[39]), .out(n1224) );
  nand2 C1839 ( .a(n1521), .b(N65), .out(n1223) );
  nand2 C1838 ( .a(n1223), .b(n1224), .out(N179) );
  nand2 C1836 ( .a(n1590), .b(final_floor_elevator1[40]), .out(n1222) );
  nand2 C1835 ( .a(n1520), .b(N66), .out(n1221) );
  nand2 C1834 ( .a(n1221), .b(n1222), .out(N178) );
  nand2 C1832 ( .a(n1590), .b(final_floor_elevator1[41]), .out(n1220) );
  nand2 C1831 ( .a(n1520), .b(N67), .out(n1219) );
  nand2 C1830 ( .a(n1219), .b(n1220), .out(N177) );
  nand2 C1828 ( .a(n1590), .b(final_floor_elevator1[42]), .out(n1218) );
  nand2 C1827 ( .a(n1520), .b(N68), .out(n1217) );
  nand2 C1826 ( .a(n1217), .b(n1218), .out(N176) );
  nand2 C1824 ( .a(n1589), .b(final_floor_elevator1[43]), .out(n1216) );
  nand2 C1823 ( .a(n1519), .b(N69), .out(n1215) );
  nand2 C1822 ( .a(n1215), .b(n1216), .out(N175) );
  nand2 C1820 ( .a(n1589), .b(final_floor_elevator1[44]), .out(n1214) );
  nand2 C1819 ( .a(n1519), .b(N70), .out(n1213) );
  nand2 C1818 ( .a(n1213), .b(n1214), .out(N174) );
  nand2 C1816 ( .a(n1589), .b(final_floor_elevator1[45]), .out(n1212) );
  nand2 C1815 ( .a(n1519), .b(N71), .out(n1211) );
  nand2 C1814 ( .a(n1211), .b(n1212), .out(N173) );
  nand2 C1812 ( .a(n1589), .b(final_floor_elevator1[46]), .out(n1210) );
  nand2 C1811 ( .a(n1518), .b(N72), .out(n1209) );
  nand2 C1810 ( .a(n1209), .b(n1210), .out(N172) );
  nand2 C1808 ( .a(n1589), .b(final_floor_elevator1[47]), .out(n1208) );
  nand2 C1807 ( .a(n1518), .b(N73), .out(n1207) );
  nand2 C1806 ( .a(n1207), .b(n1208), .out(N171) );
  nand2 C1804 ( .a(n1589), .b(final_floor_elevator1[48]), .out(n1206) );
  nand2 C1803 ( .a(n1518), .b(N74), .out(n1205) );
  nand2 C1802 ( .a(n1205), .b(n1206), .out(N170) );
  nand2 C1800 ( .a(n1589), .b(final_floor_elevator1[49]), .out(n1204) );
  nand2 C1799 ( .a(n1517), .b(N75), .out(n1203) );
  nand2 C1798 ( .a(n1203), .b(n1204), .out(N169) );
  nand2 C1796 ( .a(n1594), .b(final_floor_elevator1[50]), .out(n1202) );
  nand2 C1795 ( .a(n1513), .b(N77), .out(n1201) );
  nand2 C1794 ( .a(n1201), .b(n1202), .out(N168) );
  nand2 C1792 ( .a(n1594), .b(final_floor_elevator1[51]), .out(n1200) );
  nand2 C1791 ( .a(n1513), .b(N78), .out(n1199) );
  nand2 C1790 ( .a(n1199), .b(n1200), .out(N167) );
  nand2 C1788 ( .a(n1594), .b(final_floor_elevator1[52]), .out(n1198) );
  nand2 C1787 ( .a(n1513), .b(N79), .out(n1197) );
  nand2 C1786 ( .a(n1197), .b(n1198), .out(N166) );
  nand2 C1784 ( .a(n1594), .b(final_floor_elevator1[53]), .out(n1196) );
  nand2 C1783 ( .a(n1514), .b(N80), .out(n1195) );
  nand2 C1782 ( .a(n1195), .b(n1196), .out(N165) );
  nand2 C1780 ( .a(n1594), .b(final_floor_elevator1[54]), .out(n1194) );
  nand2 C1779 ( .a(n1514), .b(N81), .out(n1193) );
  nand2 C1778 ( .a(n1193), .b(n1194), .out(N164) );
  nand2 C1776 ( .a(n1594), .b(final_floor_elevator1[55]), .out(n1192) );
  nand2 C1775 ( .a(n1514), .b(N82), .out(n1191) );
  nand2 C1774 ( .a(n1191), .b(n1192), .out(N163) );
  nand2 C1772 ( .a(n1594), .b(final_floor_elevator1[56]), .out(n1190) );
  nand2 C1771 ( .a(n1515), .b(N83), .out(n1189) );
  nand2 C1770 ( .a(n1189), .b(n1190), .out(N162) );
  nand2 C1768 ( .a(n1594), .b(final_floor_elevator1[57]), .out(n1188) );
  nand2 C1767 ( .a(n1515), .b(N84), .out(n1187) );
  nand2 C1766 ( .a(n1187), .b(n1188), .out(N161) );
  nand2 C1764 ( .a(n1594), .b(final_floor_elevator1[58]), .out(n1186) );
  nand2 C1763 ( .a(n1515), .b(N85), .out(n1185) );
  nand2 C1762 ( .a(n1185), .b(n1186), .out(N160) );
  nand2 C1760 ( .a(n1593), .b(final_floor_elevator1[59]), .out(n1184) );
  nand2 C1759 ( .a(n1516), .b(N86), .out(n1183) );
  nand2 C1758 ( .a(n1183), .b(n1184), .out(N159) );
  nand2 C1756 ( .a(n1593), .b(final_floor_elevator1[60]), .out(n1182) );
  nand2 C1755 ( .a(n1516), .b(N87), .out(n1181) );
  nand2 C1754 ( .a(n1181), .b(n1182), .out(N158) );
  nand2 C1752 ( .a(n1593), .b(final_floor_elevator1[61]), .out(n1180) );
  nand2 C1751 ( .a(n1516), .b(N88), .out(n1179) );
  nand2 C1750 ( .a(n1179), .b(n1180), .out(N157) );
  nand2 C1748 ( .a(n1593), .b(final_floor_elevator1[62]), .out(n1178) );
  nand2 C1747 ( .a(n1517), .b(N89), .out(n1177) );
  nand2 C1746 ( .a(n1177), .b(n1178), .out(N156) );
  nand2 C1744 ( .a(n1593), .b(\ne_47/SA ), .out(n1176) );
  nand2 C1743 ( .a(n1517), .b(N90), .out(n1175) );
  nand2 C1742 ( .a(n1175), .b(n1176), .out(\r125/SA ) );
  nand2 C1740 ( .a(n1684), .b(current_floor_output_elevator1[0]), .out(n775)
         );
  nand2 C1739 ( .a(n1656), .b(current_floor_elevator1[0]), .out(n774) );
  nand2 C1736 ( .a(n1684), .b(current_floor_output_elevator1[1]), .out(n771)
         );
  nand2 C1735 ( .a(n1656), .b(current_floor_elevator1[1]), .out(n770) );
  nand2 C1732 ( .a(n1683), .b(current_floor_output_elevator1[2]), .out(n773)
         );
  nand2 C1731 ( .a(n1656), .b(current_floor_elevator1[2]), .out(n772) );
  nand2 C1728 ( .a(n1683), .b(current_floor_output_elevator1[3]), .out(n777)
         );
  nand2 C1727 ( .a(n1655), .b(current_floor_elevator1[3]), .out(n776) );
  nand2 C1724 ( .a(n1683), .b(current_floor_output_elevator1[4]), .out(n779)
         );
  nand2 C1723 ( .a(n1655), .b(current_floor_elevator1[4]), .out(n778) );
  nand2 C1720 ( .a(n1682), .b(current_floor_output_elevator1[5]), .out(n781)
         );
  nand2 C1719 ( .a(n1655), .b(current_floor_elevator1[5]), .out(n780) );
  nand2 C1716 ( .a(n1682), .b(current_floor_output_elevator1[6]), .out(n783)
         );
  nand2 C1715 ( .a(n1655), .b(current_floor_elevator1[6]), .out(n782) );
  nand2 C1712 ( .a(n1682), .b(current_floor_output_elevator1[7]), .out(n785)
         );
  nand2 C1711 ( .a(n1655), .b(current_floor_elevator1[7]), .out(n784) );
  nand2 C1708 ( .a(n1681), .b(current_floor_output_elevator1[8]), .out(n787)
         );
  nand2 C1707 ( .a(n1655), .b(current_floor_elevator1[8]), .out(n786) );
  nand2 C1704 ( .a(n1681), .b(current_floor_output_elevator1[9]), .out(n789)
         );
  nand2 C1703 ( .a(n1655), .b(current_floor_elevator1[9]), .out(n788) );
  nand2 C1700 ( .a(n1681), .b(current_floor_output_elevator1[10]), .out(n791)
         );
  nand2 C1699 ( .a(n1655), .b(current_floor_elevator1[10]), .out(n790) );
  nand2 C1696 ( .a(n1680), .b(current_floor_output_elevator1[11]), .out(n793)
         );
  nand2 C1695 ( .a(n1655), .b(current_floor_elevator1[11]), .out(n792) );
  nand2 C1692 ( .a(n1680), .b(current_floor_output_elevator1[12]), .out(n795)
         );
  nand2 C1691 ( .a(n1655), .b(current_floor_elevator1[12]), .out(n794) );
  nand2 C1688 ( .a(n1680), .b(current_floor_output_elevator1[13]), .out(n797)
         );
  nand2 C1687 ( .a(n1655), .b(current_floor_elevator1[13]), .out(n796) );
  nand2 C1684 ( .a(n1679), .b(current_floor_output_elevator1[14]), .out(n799)
         );
  nand2 C1683 ( .a(n1655), .b(current_floor_elevator1[14]), .out(n798) );
  nand2 C1680 ( .a(n1679), .b(current_floor_output_elevator1[15]), .out(n801)
         );
  nand2 C1679 ( .a(n1654), .b(current_floor_elevator1[15]), .out(n800) );
  nand2 C1676 ( .a(n1679), .b(current_floor_output_elevator1[16]), .out(n803)
         );
  nand2 C1675 ( .a(n1654), .b(current_floor_elevator1[16]), .out(n802) );
  nand2 C1672 ( .a(n1678), .b(current_floor_output_elevator1[17]), .out(n805)
         );
  nand2 C1671 ( .a(n1654), .b(current_floor_elevator1[17]), .out(n804) );
  nand2 C1668 ( .a(n1678), .b(current_floor_output_elevator1[18]), .out(n807)
         );
  nand2 C1667 ( .a(n1654), .b(current_floor_elevator1[18]), .out(n806) );
  nand2 C1664 ( .a(n1678), .b(current_floor_output_elevator1[19]), .out(n809)
         );
  nand2 C1663 ( .a(n1654), .b(current_floor_elevator1[19]), .out(n808) );
  nand2 C1660 ( .a(n1677), .b(current_floor_output_elevator1[20]), .out(n811)
         );
  nand2 C1659 ( .a(n1654), .b(current_floor_elevator1[20]), .out(n810) );
  nand2 C1656 ( .a(n1677), .b(current_floor_output_elevator1[21]), .out(n813)
         );
  nand2 C1655 ( .a(n1654), .b(current_floor_elevator1[21]), .out(n812) );
  nand2 C1652 ( .a(n1677), .b(current_floor_output_elevator1[22]), .out(n815)
         );
  nand2 C1651 ( .a(n1654), .b(current_floor_elevator1[22]), .out(n814) );
  nand2 C1648 ( .a(n1676), .b(current_floor_output_elevator1[23]), .out(n817)
         );
  nand2 C1647 ( .a(n1654), .b(current_floor_elevator1[23]), .out(n816) );
  nand2 C1644 ( .a(n1676), .b(current_floor_output_elevator1[24]), .out(n819)
         );
  nand2 C1643 ( .a(n1654), .b(current_floor_elevator1[24]), .out(n818) );
  nand2 C1640 ( .a(n1676), .b(current_floor_output_elevator1[25]), .out(n821)
         );
  nand2 C1639 ( .a(n1654), .b(current_floor_elevator1[25]), .out(n820) );
  nand2 C1636 ( .a(n1675), .b(current_floor_output_elevator1[26]), .out(n823)
         );
  nand2 C1635 ( .a(n1654), .b(current_floor_elevator1[26]), .out(n822) );
  nand2 C1632 ( .a(n1675), .b(current_floor_output_elevator1[27]), .out(n825)
         );
  nand2 C1631 ( .a(n1653), .b(current_floor_elevator1[27]), .out(n824) );
  nand2 C1628 ( .a(n1675), .b(current_floor_output_elevator1[28]), .out(n827)
         );
  nand2 C1627 ( .a(n1653), .b(current_floor_elevator1[28]), .out(n826) );
  nand2 C1624 ( .a(n1674), .b(current_floor_output_elevator1[29]), .out(n829)
         );
  nand2 C1623 ( .a(n1653), .b(current_floor_elevator1[29]), .out(n828) );
  nand2 C1620 ( .a(n1674), .b(current_floor_output_elevator1[30]), .out(n831)
         );
  nand2 C1619 ( .a(n1653), .b(current_floor_elevator1[30]), .out(n830) );
  nand2 C1616 ( .a(n1674), .b(current_floor_output_elevator1[31]), .out(n833)
         );
  nand2 C1615 ( .a(n1653), .b(current_floor_elevator1[31]), .out(n832) );
  nand2 C1612 ( .a(n1673), .b(current_floor_output_elevator1[32]), .out(n835)
         );
  nand2 C1611 ( .a(n1653), .b(current_floor_elevator1[32]), .out(n834) );
  nand2 C1608 ( .a(n1673), .b(current_floor_output_elevator1[33]), .out(n837)
         );
  nand2 C1607 ( .a(n1653), .b(current_floor_elevator1[33]), .out(n836) );
  nand2 C1604 ( .a(n1673), .b(current_floor_output_elevator1[34]), .out(n839)
         );
  nand2 C1603 ( .a(n1653), .b(current_floor_elevator1[34]), .out(n838) );
  nand2 C1600 ( .a(n1672), .b(current_floor_output_elevator1[35]), .out(n841)
         );
  nand2 C1599 ( .a(n1653), .b(current_floor_elevator1[35]), .out(n840) );
  nand2 C1596 ( .a(n1672), .b(current_floor_output_elevator1[36]), .out(n843)
         );
  nand2 C1595 ( .a(n1653), .b(current_floor_elevator1[36]), .out(n842) );
  nand2 C1592 ( .a(n1672), .b(current_floor_output_elevator1[37]), .out(n845)
         );
  nand2 C1591 ( .a(n1653), .b(current_floor_elevator1[37]), .out(n844) );
  nand2 C1588 ( .a(n1671), .b(current_floor_output_elevator1[38]), .out(n847)
         );
  nand2 C1587 ( .a(n1653), .b(current_floor_elevator1[38]), .out(n846) );
  nand2 C1584 ( .a(n1671), .b(current_floor_output_elevator1[39]), .out(n849)
         );
  nand2 C1583 ( .a(n1652), .b(current_floor_elevator1[39]), .out(n848) );
  nand2 C1580 ( .a(n1671), .b(current_floor_output_elevator1[40]), .out(n851)
         );
  nand2 C1579 ( .a(n1652), .b(current_floor_elevator1[40]), .out(n850) );
  nand2 C1576 ( .a(n1670), .b(current_floor_output_elevator1[41]), .out(n853)
         );
  nand2 C1575 ( .a(n1652), .b(current_floor_elevator1[41]), .out(n852) );
  nand2 C1572 ( .a(n1670), .b(current_floor_output_elevator1[42]), .out(n855)
         );
  nand2 C1571 ( .a(n1652), .b(current_floor_elevator1[42]), .out(n854) );
  nand2 C1568 ( .a(n1670), .b(current_floor_output_elevator1[43]), .out(n857)
         );
  nand2 C1567 ( .a(n1652), .b(current_floor_elevator1[43]), .out(n856) );
  nand2 C1564 ( .a(n1669), .b(current_floor_output_elevator1[44]), .out(n859)
         );
  nand2 C1563 ( .a(n1652), .b(current_floor_elevator1[44]), .out(n858) );
  nand2 C1560 ( .a(n1669), .b(current_floor_output_elevator1[45]), .out(n861)
         );
  nand2 C1559 ( .a(n1652), .b(current_floor_elevator1[45]), .out(n860) );
  nand2 C1556 ( .a(n1669), .b(current_floor_output_elevator1[46]), .out(n863)
         );
  nand2 C1555 ( .a(n1652), .b(current_floor_elevator1[46]), .out(n862) );
  nand2 C1552 ( .a(n1668), .b(current_floor_output_elevator1[47]), .out(n865)
         );
  nand2 C1551 ( .a(n1652), .b(current_floor_elevator1[47]), .out(n864) );
  nand2 C1548 ( .a(n1668), .b(current_floor_output_elevator1[48]), .out(n867)
         );
  nand2 C1547 ( .a(n1652), .b(current_floor_elevator1[48]), .out(n866) );
  nand2 C1544 ( .a(n1668), .b(current_floor_output_elevator1[49]), .out(n869)
         );
  nand2 C1543 ( .a(n1652), .b(current_floor_elevator1[49]), .out(n868) );
  nand2 C1540 ( .a(n1667), .b(current_floor_output_elevator1[50]), .out(n871)
         );
  nand2 C1539 ( .a(n1652), .b(current_floor_elevator1[50]), .out(n870) );
  nand2 C1536 ( .a(n1667), .b(current_floor_output_elevator1[51]), .out(n873)
         );
  nand2 C1535 ( .a(n1651), .b(current_floor_elevator1[51]), .out(n872) );
  nand2 C1532 ( .a(n1667), .b(current_floor_output_elevator1[52]), .out(n875)
         );
  nand2 C1531 ( .a(n1651), .b(current_floor_elevator1[52]), .out(n874) );
  nand2 C1528 ( .a(n1666), .b(current_floor_output_elevator1[53]), .out(n877)
         );
  nand2 C1527 ( .a(n1651), .b(current_floor_elevator1[53]), .out(n876) );
  nand2 C1524 ( .a(n1666), .b(current_floor_output_elevator1[54]), .out(n879)
         );
  nand2 C1523 ( .a(n1651), .b(current_floor_elevator1[54]), .out(n878) );
  nand2 C1520 ( .a(n1666), .b(current_floor_output_elevator1[55]), .out(n881)
         );
  nand2 C1519 ( .a(n1651), .b(current_floor_elevator1[55]), .out(n880) );
  nand2 C1516 ( .a(n1665), .b(current_floor_output_elevator1[56]), .out(n883)
         );
  nand2 C1515 ( .a(n1651), .b(current_floor_elevator1[56]), .out(n882) );
  nand2 C1512 ( .a(n1665), .b(current_floor_output_elevator1[57]), .out(n885)
         );
  nand2 C1511 ( .a(n1651), .b(current_floor_elevator1[57]), .out(n884) );
  nand2 C1508 ( .a(n1665), .b(current_floor_output_elevator1[58]), .out(n887)
         );
  nand2 C1507 ( .a(n1651), .b(current_floor_elevator1[58]), .out(n886) );
  nand2 C1504 ( .a(n1664), .b(current_floor_output_elevator1[59]), .out(n889)
         );
  nand2 C1503 ( .a(n1651), .b(current_floor_elevator1[59]), .out(n888) );
  nand2 C1500 ( .a(n1664), .b(current_floor_output_elevator1[60]), .out(n891)
         );
  nand2 C1499 ( .a(n1651), .b(current_floor_elevator1[60]), .out(n890) );
  nand2 C1496 ( .a(n1664), .b(current_floor_output_elevator1[61]), .out(n893)
         );
  nand2 C1495 ( .a(n1651), .b(current_floor_elevator1[61]), .out(n892) );
  nand2 C1492 ( .a(n1663), .b(current_floor_output_elevator1[62]), .out(n895)
         );
  nand2 C1491 ( .a(n1651), .b(current_floor_elevator1[62]), .out(n894) );
  nand2 C1488 ( .a(n1663), .b(\eq_42_3/SA ), .out(n897) );
  nand2 C1487 ( .a(n1650), .b(current_floor_elevator1[63]), .out(n896) );
  nand2 C1478 ( .a(N604), .b(N605), .out(n1174) );
  nand2 C1477 ( .a(N609), .b(N15), .out(n640) );
  nand2 C1475 ( .a(N606), .b(N605), .out(n1173) );
  nand2 C1474 ( .a(N607), .b(N12), .out(n641) );
  inv I_4 ( .in(elevator1_status), .out(N606) );
  inv I_3 ( .in(request_taken), .out(N605) );
  inv I_2 ( .in(elevator2_status), .out(N604) );
  dff emergency_signal_elevator2_reg ( .d(N514), .gclk(clk), .rnot(1'b1), .q(
        emergency_signal_elevator2) );
  dff emergency_signal_elevator1_reg ( .d(N230), .gclk(clk), .rnot(1'b1), .q(
        emergency_signal_elevator1) );
  dff request_taken_reg ( .d(n1162), .gclk(clk), .rnot(1'b1), .q(request_taken) );
  dff \final_floor_elevator1_reg[50]  ( .d(n1161), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator1[50]) );
  dff \final_floor_elevator1_reg[51]  ( .d(n1160), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator1[51]) );
  dff \final_floor_elevator1_reg[52]  ( .d(n1159), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator1[52]) );
  dff \final_floor_elevator1_reg[53]  ( .d(n1158), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator1[53]) );
  dff \final_floor_elevator1_reg[54]  ( .d(n1157), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator1[54]) );
  dff \final_floor_elevator1_reg[55]  ( .d(n1156), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator1[55]) );
  dff \final_floor_elevator1_reg[56]  ( .d(n1155), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator1[56]) );
  dff \final_floor_elevator1_reg[57]  ( .d(n1154), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator1[57]) );
  dff \final_floor_elevator1_reg[58]  ( .d(n1153), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator1[58]) );
  dff \final_floor_elevator1_reg[59]  ( .d(n1152), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator1[59]) );
  dff \final_floor_elevator1_reg[60]  ( .d(n1151), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator1[60]) );
  dff \final_floor_elevator1_reg[61]  ( .d(n1150), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator1[61]) );
  dff \final_floor_elevator1_reg[62]  ( .d(n1149), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator1[62]) );
  dff \final_floor_elevator1_reg[63]  ( .d(n1148), .gclk(clk), .rnot(1'b1), 
        .q(\ne_47/SA ) );
  dff \final_floor_elevator1_reg[49]  ( .d(n1147), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator1[49]) );
  dff \final_floor_elevator1_reg[48]  ( .d(n1146), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator1[48]) );
  dff \final_floor_elevator1_reg[47]  ( .d(n1145), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator1[47]) );
  dff \final_floor_elevator1_reg[46]  ( .d(n1144), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator1[46]) );
  dff \final_floor_elevator1_reg[45]  ( .d(n1143), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator1[45]) );
  dff \final_floor_elevator1_reg[44]  ( .d(n1142), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator1[44]) );
  dff \final_floor_elevator1_reg[43]  ( .d(n1141), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator1[43]) );
  dff \final_floor_elevator1_reg[42]  ( .d(n1140), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator1[42]) );
  dff \final_floor_elevator1_reg[41]  ( .d(n1139), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator1[41]) );
  dff \final_floor_elevator1_reg[40]  ( .d(n1138), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator1[40]) );
  dff \final_floor_elevator1_reg[39]  ( .d(n1137), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator1[39]) );
  dff \final_floor_elevator1_reg[38]  ( .d(n1136), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator1[38]) );
  dff \final_floor_elevator1_reg[37]  ( .d(n1135), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator1[37]) );
  dff \final_floor_elevator1_reg[36]  ( .d(n1134), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator1[36]) );
  dff \final_floor_elevator1_reg[35]  ( .d(n1133), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator1[35]) );
  dff \final_floor_elevator1_reg[34]  ( .d(n1132), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator1[34]) );
  dff \final_floor_elevator1_reg[33]  ( .d(n1131), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator1[33]) );
  dff \final_floor_elevator1_reg[32]  ( .d(n1130), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator1[32]) );
  dff \final_floor_elevator1_reg[31]  ( .d(n1129), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator1[31]) );
  dff \final_floor_elevator1_reg[30]  ( .d(n1128), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator1[30]) );
  dff \final_floor_elevator1_reg[29]  ( .d(n1127), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator1[29]) );
  dff \final_floor_elevator1_reg[28]  ( .d(n1126), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator1[28]) );
  dff \final_floor_elevator1_reg[27]  ( .d(n1125), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator1[27]) );
  dff \final_floor_elevator1_reg[26]  ( .d(n1124), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator1[26]) );
  dff \final_floor_elevator1_reg[25]  ( .d(n1123), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator1[25]) );
  dff \final_floor_elevator1_reg[24]  ( .d(n1122), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator1[24]) );
  dff \final_floor_elevator1_reg[23]  ( .d(n1121), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator1[23]) );
  dff \final_floor_elevator1_reg[22]  ( .d(n1120), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator1[22]) );
  dff \final_floor_elevator1_reg[21]  ( .d(n1119), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator1[21]) );
  dff \final_floor_elevator1_reg[20]  ( .d(n1118), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator1[20]) );
  dff \final_floor_elevator1_reg[19]  ( .d(n1117), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator1[19]) );
  dff \final_floor_elevator1_reg[18]  ( .d(n1116), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator1[18]) );
  dff \final_floor_elevator1_reg[17]  ( .d(n1115), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator1[17]) );
  dff \final_floor_elevator1_reg[16]  ( .d(n1114), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator1[16]) );
  dff \final_floor_elevator1_reg[15]  ( .d(n1113), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator1[15]) );
  dff \final_floor_elevator1_reg[14]  ( .d(n1112), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator1[14]) );
  dff \final_floor_elevator1_reg[13]  ( .d(n1111), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator1[13]) );
  dff \final_floor_elevator1_reg[12]  ( .d(n1110), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator1[12]) );
  dff \final_floor_elevator1_reg[11]  ( .d(n1109), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator1[11]) );
  dff \final_floor_elevator1_reg[10]  ( .d(n1108), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator1[10]) );
  dff \final_floor_elevator1_reg[9]  ( .d(n1107), .gclk(clk), .rnot(1'b1), .q(
        final_floor_elevator1[9]) );
  dff \final_floor_elevator1_reg[8]  ( .d(n1106), .gclk(clk), .rnot(1'b1), .q(
        final_floor_elevator1[8]) );
  dff \final_floor_elevator1_reg[7]  ( .d(n1105), .gclk(clk), .rnot(1'b1), .q(
        final_floor_elevator1[7]) );
  dff \final_floor_elevator1_reg[6]  ( .d(n1104), .gclk(clk), .rnot(1'b1), .q(
        final_floor_elevator1[6]) );
  dff \final_floor_elevator1_reg[5]  ( .d(n1103), .gclk(clk), .rnot(1'b1), .q(
        final_floor_elevator1[5]) );
  dff \final_floor_elevator1_reg[4]  ( .d(n1102), .gclk(clk), .rnot(1'b1), .q(
        final_floor_elevator1[4]) );
  dff \final_floor_elevator1_reg[3]  ( .d(n1101), .gclk(clk), .rnot(1'b1), .q(
        final_floor_elevator1[3]) );
  dff \final_floor_elevator1_reg[2]  ( .d(n1100), .gclk(clk), .rnot(1'b1), .q(
        final_floor_elevator1[2]) );
  dff \final_floor_elevator1_reg[1]  ( .d(n1099), .gclk(clk), .rnot(1'b1), .q(
        final_floor_elevator1[1]) );
  dff \final_floor_elevator1_reg[0]  ( .d(n1098), .gclk(clk), .rnot(1'b1), .q(
        final_floor_elevator1[0]) );
  dff \final_floor_elevator2_reg[50]  ( .d(n1097), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator2[50]) );
  dff \final_floor_elevator2_reg[51]  ( .d(n1096), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator2[51]) );
  dff \final_floor_elevator2_reg[52]  ( .d(n1095), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator2[52]) );
  dff \final_floor_elevator2_reg[53]  ( .d(n1094), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator2[53]) );
  dff \final_floor_elevator2_reg[54]  ( .d(n1093), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator2[54]) );
  dff \final_floor_elevator2_reg[55]  ( .d(n1092), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator2[55]) );
  dff \final_floor_elevator2_reg[56]  ( .d(n1091), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator2[56]) );
  dff \final_floor_elevator2_reg[57]  ( .d(n1090), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator2[57]) );
  dff \final_floor_elevator2_reg[58]  ( .d(n1089), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator2[58]) );
  dff \final_floor_elevator2_reg[59]  ( .d(n1088), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator2[59]) );
  dff \final_floor_elevator2_reg[60]  ( .d(n1087), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator2[60]) );
  dff \final_floor_elevator2_reg[61]  ( .d(n1086), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator2[61]) );
  dff \final_floor_elevator2_reg[62]  ( .d(n1085), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator2[62]) );
  dff \final_floor_elevator2_reg[63]  ( .d(n1084), .gclk(clk), .rnot(1'b1), 
        .q(\ne_42/SA ) );
  dff \final_floor_elevator2_reg[49]  ( .d(n1083), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator2[49]) );
  dff \final_floor_elevator2_reg[48]  ( .d(n1082), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator2[48]) );
  dff \final_floor_elevator2_reg[47]  ( .d(n1081), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator2[47]) );
  dff \final_floor_elevator2_reg[46]  ( .d(n1080), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator2[46]) );
  dff \final_floor_elevator2_reg[45]  ( .d(n1079), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator2[45]) );
  dff \final_floor_elevator2_reg[44]  ( .d(n1078), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator2[44]) );
  dff \final_floor_elevator2_reg[43]  ( .d(n1077), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator2[43]) );
  dff \final_floor_elevator2_reg[42]  ( .d(n1076), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator2[42]) );
  dff \final_floor_elevator2_reg[41]  ( .d(n1075), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator2[41]) );
  dff \final_floor_elevator2_reg[40]  ( .d(n1074), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator2[40]) );
  dff \final_floor_elevator2_reg[39]  ( .d(n1073), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator2[39]) );
  dff \final_floor_elevator2_reg[38]  ( .d(n1072), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator2[38]) );
  dff \final_floor_elevator2_reg[37]  ( .d(n1071), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator2[37]) );
  dff \final_floor_elevator2_reg[36]  ( .d(n1070), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator2[36]) );
  dff \final_floor_elevator2_reg[35]  ( .d(n1069), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator2[35]) );
  dff \final_floor_elevator2_reg[34]  ( .d(n1068), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator2[34]) );
  dff \final_floor_elevator2_reg[33]  ( .d(n1067), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator2[33]) );
  dff \final_floor_elevator2_reg[32]  ( .d(n1066), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator2[32]) );
  dff \final_floor_elevator2_reg[31]  ( .d(n1065), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator2[31]) );
  dff \final_floor_elevator2_reg[30]  ( .d(n1064), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator2[30]) );
  dff \final_floor_elevator2_reg[29]  ( .d(n1063), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator2[29]) );
  dff \final_floor_elevator2_reg[28]  ( .d(n1062), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator2[28]) );
  dff \final_floor_elevator2_reg[27]  ( .d(n1061), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator2[27]) );
  dff \final_floor_elevator2_reg[26]  ( .d(n1060), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator2[26]) );
  dff \final_floor_elevator2_reg[25]  ( .d(n1059), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator2[25]) );
  dff \final_floor_elevator2_reg[24]  ( .d(n1058), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator2[24]) );
  dff \final_floor_elevator2_reg[23]  ( .d(n1057), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator2[23]) );
  dff \final_floor_elevator2_reg[22]  ( .d(n1056), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator2[22]) );
  dff \final_floor_elevator2_reg[21]  ( .d(n1055), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator2[21]) );
  dff \final_floor_elevator2_reg[20]  ( .d(n1054), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator2[20]) );
  dff \final_floor_elevator2_reg[19]  ( .d(n1053), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator2[19]) );
  dff \final_floor_elevator2_reg[18]  ( .d(n1052), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator2[18]) );
  dff \final_floor_elevator2_reg[17]  ( .d(n1051), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator2[17]) );
  dff \final_floor_elevator2_reg[16]  ( .d(n1050), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator2[16]) );
  dff \final_floor_elevator2_reg[15]  ( .d(n1049), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator2[15]) );
  dff \final_floor_elevator2_reg[14]  ( .d(n1048), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator2[14]) );
  dff \final_floor_elevator2_reg[13]  ( .d(n1047), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator2[13]) );
  dff \final_floor_elevator2_reg[12]  ( .d(n1046), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator2[12]) );
  dff \final_floor_elevator2_reg[11]  ( .d(n1045), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator2[11]) );
  dff \final_floor_elevator2_reg[10]  ( .d(n1044), .gclk(clk), .rnot(1'b1), 
        .q(final_floor_elevator2[10]) );
  dff \final_floor_elevator2_reg[9]  ( .d(n1043), .gclk(clk), .rnot(1'b1), .q(
        final_floor_elevator2[9]) );
  dff \final_floor_elevator2_reg[8]  ( .d(n1042), .gclk(clk), .rnot(1'b1), .q(
        final_floor_elevator2[8]) );
  dff \final_floor_elevator2_reg[7]  ( .d(n1041), .gclk(clk), .rnot(1'b1), .q(
        final_floor_elevator2[7]) );
  dff \final_floor_elevator2_reg[6]  ( .d(n1040), .gclk(clk), .rnot(1'b1), .q(
        final_floor_elevator2[6]) );
  dff \final_floor_elevator2_reg[5]  ( .d(n1039), .gclk(clk), .rnot(1'b1), .q(
        final_floor_elevator2[5]) );
  dff \final_floor_elevator2_reg[4]  ( .d(n1038), .gclk(clk), .rnot(1'b1), .q(
        final_floor_elevator2[4]) );
  dff \final_floor_elevator2_reg[3]  ( .d(n1037), .gclk(clk), .rnot(1'b1), .q(
        final_floor_elevator2[3]) );
  dff \final_floor_elevator2_reg[2]  ( .d(n1036), .gclk(clk), .rnot(1'b1), .q(
        final_floor_elevator2[2]) );
  dff \final_floor_elevator2_reg[1]  ( .d(n1035), .gclk(clk), .rnot(1'b1), .q(
        final_floor_elevator2[1]) );
  dff \final_floor_elevator2_reg[0]  ( .d(n1034), .gclk(clk), .rnot(1'b1), .q(
        final_floor_elevator2[0]) );
  dff \current_floor_output_elevator2_reg[0]  ( .d(n1033), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator2[0]) );
  dff \current_floor_output_elevator2_reg[1]  ( .d(n1032), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator2[1]) );
  dff \current_floor_output_elevator2_reg[2]  ( .d(n1031), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator2[2]) );
  dff \current_floor_output_elevator2_reg[3]  ( .d(n1030), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator2[3]) );
  dff \current_floor_output_elevator2_reg[4]  ( .d(n1029), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator2[4]) );
  dff \current_floor_output_elevator2_reg[5]  ( .d(n1028), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator2[5]) );
  dff \current_floor_output_elevator2_reg[6]  ( .d(n1027), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator2[6]) );
  dff \current_floor_output_elevator2_reg[7]  ( .d(n1026), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator2[7]) );
  dff \current_floor_output_elevator2_reg[8]  ( .d(n1025), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator2[8]) );
  dff \current_floor_output_elevator2_reg[9]  ( .d(n1024), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator2[9]) );
  dff \current_floor_output_elevator2_reg[10]  ( .d(n1023), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator2[10]) );
  dff \current_floor_output_elevator2_reg[11]  ( .d(n1022), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator2[11]) );
  dff \current_floor_output_elevator2_reg[12]  ( .d(n1021), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator2[12]) );
  dff \current_floor_output_elevator2_reg[13]  ( .d(n1020), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator2[13]) );
  dff \current_floor_output_elevator2_reg[14]  ( .d(n1019), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator2[14]) );
  dff \current_floor_output_elevator2_reg[15]  ( .d(n1018), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator2[15]) );
  dff \current_floor_output_elevator2_reg[16]  ( .d(n1017), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator2[16]) );
  dff \current_floor_output_elevator2_reg[17]  ( .d(n1016), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator2[17]) );
  dff \current_floor_output_elevator2_reg[18]  ( .d(n1015), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator2[18]) );
  dff \current_floor_output_elevator2_reg[19]  ( .d(n1014), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator2[19]) );
  dff \current_floor_output_elevator2_reg[20]  ( .d(n1013), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator2[20]) );
  dff \current_floor_output_elevator2_reg[21]  ( .d(n1012), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator2[21]) );
  dff \current_floor_output_elevator2_reg[22]  ( .d(n1011), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator2[22]) );
  dff \current_floor_output_elevator2_reg[23]  ( .d(n1010), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator2[23]) );
  dff \current_floor_output_elevator2_reg[24]  ( .d(n1009), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator2[24]) );
  dff \current_floor_output_elevator2_reg[25]  ( .d(n1008), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator2[25]) );
  dff \current_floor_output_elevator2_reg[26]  ( .d(n1007), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator2[26]) );
  dff \current_floor_output_elevator2_reg[27]  ( .d(n1006), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator2[27]) );
  dff \current_floor_output_elevator2_reg[28]  ( .d(n1005), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator2[28]) );
  dff \current_floor_output_elevator2_reg[29]  ( .d(n1004), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator2[29]) );
  dff \current_floor_output_elevator2_reg[30]  ( .d(n1003), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator2[30]) );
  dff \current_floor_output_elevator2_reg[31]  ( .d(n1002), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator2[31]) );
  dff \current_floor_output_elevator2_reg[32]  ( .d(n1001), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator2[32]) );
  dff \current_floor_output_elevator2_reg[33]  ( .d(n1000), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator2[33]) );
  dff \current_floor_output_elevator2_reg[34]  ( .d(n999), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator2[34]) );
  dff \current_floor_output_elevator2_reg[35]  ( .d(n998), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator2[35]) );
  dff \current_floor_output_elevator2_reg[36]  ( .d(n997), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator2[36]) );
  dff \current_floor_output_elevator2_reg[37]  ( .d(n996), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator2[37]) );
  dff \current_floor_output_elevator2_reg[38]  ( .d(n995), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator2[38]) );
  dff \current_floor_output_elevator2_reg[39]  ( .d(n994), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator2[39]) );
  dff \current_floor_output_elevator2_reg[40]  ( .d(n993), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator2[40]) );
  dff \current_floor_output_elevator2_reg[41]  ( .d(n992), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator2[41]) );
  dff \current_floor_output_elevator2_reg[42]  ( .d(n991), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator2[42]) );
  dff \current_floor_output_elevator2_reg[43]  ( .d(n990), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator2[43]) );
  dff \current_floor_output_elevator2_reg[44]  ( .d(n989), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator2[44]) );
  dff \current_floor_output_elevator2_reg[45]  ( .d(n988), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator2[45]) );
  dff \current_floor_output_elevator2_reg[46]  ( .d(n987), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator2[46]) );
  dff \current_floor_output_elevator2_reg[47]  ( .d(n986), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator2[47]) );
  dff \current_floor_output_elevator2_reg[48]  ( .d(n985), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator2[48]) );
  dff \current_floor_output_elevator2_reg[49]  ( .d(n984), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator2[49]) );
  dff \current_floor_output_elevator2_reg[50]  ( .d(n983), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator2[50]) );
  dff \current_floor_output_elevator2_reg[51]  ( .d(n982), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator2[51]) );
  dff \current_floor_output_elevator2_reg[52]  ( .d(n981), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator2[52]) );
  dff \current_floor_output_elevator2_reg[53]  ( .d(n980), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator2[53]) );
  dff \current_floor_output_elevator2_reg[54]  ( .d(n979), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator2[54]) );
  dff \current_floor_output_elevator2_reg[55]  ( .d(n978), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator2[55]) );
  dff \current_floor_output_elevator2_reg[56]  ( .d(n977), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator2[56]) );
  dff \current_floor_output_elevator2_reg[57]  ( .d(n976), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator2[57]) );
  dff \current_floor_output_elevator2_reg[58]  ( .d(n975), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator2[58]) );
  dff \current_floor_output_elevator2_reg[59]  ( .d(n974), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator2[59]) );
  dff \current_floor_output_elevator2_reg[60]  ( .d(n973), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator2[60]) );
  dff \current_floor_output_elevator2_reg[61]  ( .d(n972), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator2[61]) );
  dff \current_floor_output_elevator2_reg[62]  ( .d(n971), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator2[62]) );
  dff \current_floor_output_elevator2_reg[63]  ( .d(n970), .gclk(clk), .rnot(
        1'b1), .q(\eq_47_3/SA ) );
  dff elevator2_status_reg ( .d(n969), .gclk(clk), .rnot(1'b1), .q(
        elevator2_status) );
  dff \direction_elevator2_reg[1]  ( .d(n968), .gclk(clk), .rnot(1'b1), .q(
        direction_elevator2[1]) );
  dff arrived_elevator2_reg ( .d(n967), .gclk(clk), .rnot(1'b1), .q(
        arrived_elevator2) );
  dff \direction_elevator2_reg[0]  ( .d(n966), .gclk(clk), .rnot(1'b1), .q(
        direction_elevator2[0]) );
  dff \current_floor_output_elevator1_reg[0]  ( .d(n965), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator1[0]) );
  dff \current_floor_output_elevator1_reg[1]  ( .d(n964), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator1[1]) );
  dff \current_floor_output_elevator1_reg[2]  ( .d(n963), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator1[2]) );
  dff \current_floor_output_elevator1_reg[3]  ( .d(n962), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator1[3]) );
  dff \current_floor_output_elevator1_reg[4]  ( .d(n961), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator1[4]) );
  dff \current_floor_output_elevator1_reg[5]  ( .d(n960), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator1[5]) );
  dff \current_floor_output_elevator1_reg[6]  ( .d(n959), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator1[6]) );
  dff \current_floor_output_elevator1_reg[7]  ( .d(n958), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator1[7]) );
  dff \current_floor_output_elevator1_reg[8]  ( .d(n957), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator1[8]) );
  dff \current_floor_output_elevator1_reg[9]  ( .d(n956), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator1[9]) );
  dff \current_floor_output_elevator1_reg[10]  ( .d(n955), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator1[10]) );
  dff \current_floor_output_elevator1_reg[11]  ( .d(n954), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator1[11]) );
  dff \current_floor_output_elevator1_reg[12]  ( .d(n953), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator1[12]) );
  dff \current_floor_output_elevator1_reg[13]  ( .d(n952), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator1[13]) );
  dff \current_floor_output_elevator1_reg[14]  ( .d(n951), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator1[14]) );
  dff \current_floor_output_elevator1_reg[15]  ( .d(n950), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator1[15]) );
  dff \current_floor_output_elevator1_reg[16]  ( .d(n949), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator1[16]) );
  dff \current_floor_output_elevator1_reg[17]  ( .d(n948), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator1[17]) );
  dff \current_floor_output_elevator1_reg[18]  ( .d(n947), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator1[18]) );
  dff \current_floor_output_elevator1_reg[19]  ( .d(n946), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator1[19]) );
  dff \current_floor_output_elevator1_reg[20]  ( .d(n945), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator1[20]) );
  dff \current_floor_output_elevator1_reg[21]  ( .d(n944), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator1[21]) );
  dff \current_floor_output_elevator1_reg[22]  ( .d(n943), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator1[22]) );
  dff \current_floor_output_elevator1_reg[23]  ( .d(n942), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator1[23]) );
  dff \current_floor_output_elevator1_reg[24]  ( .d(n941), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator1[24]) );
  dff \current_floor_output_elevator1_reg[25]  ( .d(n940), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator1[25]) );
  dff \current_floor_output_elevator1_reg[26]  ( .d(n939), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator1[26]) );
  dff \current_floor_output_elevator1_reg[27]  ( .d(n938), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator1[27]) );
  dff \current_floor_output_elevator1_reg[28]  ( .d(n937), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator1[28]) );
  dff \current_floor_output_elevator1_reg[29]  ( .d(n936), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator1[29]) );
  dff \current_floor_output_elevator1_reg[30]  ( .d(n935), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator1[30]) );
  dff \current_floor_output_elevator1_reg[31]  ( .d(n934), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator1[31]) );
  dff \current_floor_output_elevator1_reg[32]  ( .d(n933), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator1[32]) );
  dff \current_floor_output_elevator1_reg[33]  ( .d(n932), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator1[33]) );
  dff \current_floor_output_elevator1_reg[34]  ( .d(n931), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator1[34]) );
  dff \current_floor_output_elevator1_reg[35]  ( .d(n930), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator1[35]) );
  dff \current_floor_output_elevator1_reg[36]  ( .d(n929), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator1[36]) );
  dff \current_floor_output_elevator1_reg[37]  ( .d(n928), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator1[37]) );
  dff \current_floor_output_elevator1_reg[38]  ( .d(n927), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator1[38]) );
  dff \current_floor_output_elevator1_reg[39]  ( .d(n926), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator1[39]) );
  dff \current_floor_output_elevator1_reg[40]  ( .d(n925), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator1[40]) );
  dff \current_floor_output_elevator1_reg[41]  ( .d(n924), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator1[41]) );
  dff \current_floor_output_elevator1_reg[42]  ( .d(n923), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator1[42]) );
  dff \current_floor_output_elevator1_reg[43]  ( .d(n922), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator1[43]) );
  dff \current_floor_output_elevator1_reg[44]  ( .d(n921), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator1[44]) );
  dff \current_floor_output_elevator1_reg[45]  ( .d(n920), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator1[45]) );
  dff \current_floor_output_elevator1_reg[46]  ( .d(n919), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator1[46]) );
  dff \current_floor_output_elevator1_reg[47]  ( .d(n918), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator1[47]) );
  dff \current_floor_output_elevator1_reg[48]  ( .d(n917), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator1[48]) );
  dff \current_floor_output_elevator1_reg[49]  ( .d(n916), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator1[49]) );
  dff \current_floor_output_elevator1_reg[50]  ( .d(n915), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator1[50]) );
  dff \current_floor_output_elevator1_reg[51]  ( .d(n914), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator1[51]) );
  dff \current_floor_output_elevator1_reg[52]  ( .d(n913), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator1[52]) );
  dff \current_floor_output_elevator1_reg[53]  ( .d(n912), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator1[53]) );
  dff \current_floor_output_elevator1_reg[54]  ( .d(n911), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator1[54]) );
  dff \current_floor_output_elevator1_reg[55]  ( .d(n910), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator1[55]) );
  dff \current_floor_output_elevator1_reg[56]  ( .d(n909), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator1[56]) );
  dff \current_floor_output_elevator1_reg[57]  ( .d(n908), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator1[57]) );
  dff \current_floor_output_elevator1_reg[58]  ( .d(n907), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator1[58]) );
  dff \current_floor_output_elevator1_reg[59]  ( .d(n906), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator1[59]) );
  dff \current_floor_output_elevator1_reg[60]  ( .d(n905), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator1[60]) );
  dff \current_floor_output_elevator1_reg[61]  ( .d(n904), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator1[61]) );
  dff \current_floor_output_elevator1_reg[62]  ( .d(n903), .gclk(clk), .rnot(
        1'b1), .q(current_floor_output_elevator1[62]) );
  dff \current_floor_output_elevator1_reg[63]  ( .d(n902), .gclk(clk), .rnot(
        1'b1), .q(\eq_42_3/SA ) );
  dff elevator1_status_reg ( .d(n901), .gclk(clk), .rnot(1'b1), .q(
        elevator1_status) );
  dff \direction_elevator1_reg[1]  ( .d(n900), .gclk(clk), .rnot(1'b1), .q(
        direction_elevator1[1]) );
  dff arrived_elevator1_reg ( .d(n899), .gclk(clk), .rnot(1'b1), .q(
        arrived_elevator1) );
  dff \direction_elevator1_reg[0]  ( .d(n898), .gclk(clk), .rnot(1'b1), .q(
        direction_elevator1[0]) );
  oai12 U3 ( .b(n18), .c(N605), .a(n19), .out(n1162) );
  nand4 U10 ( .a(n20), .b(n21), .c(n22), .d(n18), .out(n19) );
  nor2 U11 ( .a(n1595), .b(n1640), .out(n22) );
  nand3 U12 ( .a(n23), .b(n1166), .c(n24), .out(n21) );
  inv U13 ( .in(n25), .out(n24) );
  nor2 U14 ( .a(n1172), .b(N225), .out(n25) );
  nand3 U15 ( .a(n26), .b(n1168), .c(n27), .out(n20) );
  nand2 U16 ( .a(n28), .b(n29), .out(n27) );
  inv U17 ( .in(N509), .out(n29) );
  nand4 U18 ( .a(n1589), .b(n1618), .c(n32), .d(n33), .out(n18) );
  aoi12 U19 ( .b(N16), .c(n34), .a(n35), .out(n33) );
  inv U20 ( .in(n36), .out(n1043) );
  aoi22 U21 ( .a(n1507), .b(final_floor_elevator2[9]), .c(n1473), .d(N319), 
        .out(n36) );
  inv U22 ( .in(n38), .out(n1042) );
  aoi22 U23 ( .a(n1507), .b(final_floor_elevator2[8]), .c(n1473), .d(N318), 
        .out(n38) );
  inv U24 ( .in(n39), .out(n1041) );
  aoi22 U25 ( .a(n1507), .b(final_floor_elevator2[7]), .c(n1472), .d(N317), 
        .out(n39) );
  inv U26 ( .in(n40), .out(n1040) );
  aoi22 U27 ( .a(n1507), .b(final_floor_elevator2[6]), .c(n1472), .d(N316), 
        .out(n40) );
  inv U28 ( .in(n41), .out(n1084) );
  aoi22 U29 ( .a(n1472), .b(N374), .c(n1506), .d(\ne_42/SA ), .out(n41) );
  inv U30 ( .in(n42), .out(n1085) );
  aoi22 U31 ( .a(n1471), .b(N373), .c(n1506), .d(final_floor_elevator2[62]), 
        .out(n42) );
  inv U32 ( .in(n43), .out(n1086) );
  aoi22 U33 ( .a(n1471), .b(N372), .c(n1506), .d(final_floor_elevator2[61]), 
        .out(n43) );
  inv U34 ( .in(n44), .out(n1087) );
  aoi22 U35 ( .a(n1471), .b(N371), .c(n1506), .d(final_floor_elevator2[60]), 
        .out(n44) );
  inv U36 ( .in(n45), .out(n1039) );
  aoi22 U37 ( .a(n1506), .b(final_floor_elevator2[5]), .c(n1470), .d(N315), 
        .out(n45) );
  inv U38 ( .in(n46), .out(n1088) );
  aoi22 U39 ( .a(n1470), .b(N370), .c(n1506), .d(final_floor_elevator2[59]), 
        .out(n46) );
  inv U40 ( .in(n47), .out(n1089) );
  aoi22 U41 ( .a(n1470), .b(N369), .c(n1506), .d(final_floor_elevator2[58]), 
        .out(n47) );
  inv U42 ( .in(n48), .out(n1090) );
  aoi22 U43 ( .a(n1469), .b(N368), .c(n1506), .d(final_floor_elevator2[57]), 
        .out(n48) );
  inv U44 ( .in(n49), .out(n1091) );
  aoi22 U45 ( .a(n1469), .b(N367), .c(n1506), .d(final_floor_elevator2[56]), 
        .out(n49) );
  inv U46 ( .in(n50), .out(n1092) );
  aoi22 U47 ( .a(n1469), .b(N366), .c(n1506), .d(final_floor_elevator2[55]), 
        .out(n50) );
  inv U48 ( .in(n51), .out(n1093) );
  aoi22 U49 ( .a(n1468), .b(N365), .c(n1506), .d(final_floor_elevator2[54]), 
        .out(n51) );
  inv U50 ( .in(n52), .out(n1094) );
  aoi22 U51 ( .a(n1468), .b(N364), .c(n1506), .d(final_floor_elevator2[53]), 
        .out(n52) );
  inv U52 ( .in(n53), .out(n1095) );
  aoi22 U53 ( .a(n1468), .b(N363), .c(n1505), .d(final_floor_elevator2[52]), 
        .out(n53) );
  inv U54 ( .in(n54), .out(n1096) );
  aoi22 U55 ( .a(n1467), .b(N362), .c(n1505), .d(final_floor_elevator2[51]), 
        .out(n54) );
  inv U56 ( .in(n55), .out(n1097) );
  aoi22 U57 ( .a(n1467), .b(N361), .c(n1505), .d(final_floor_elevator2[50]), 
        .out(n55) );
  inv U58 ( .in(n56), .out(n1038) );
  aoi22 U59 ( .a(n1505), .b(final_floor_elevator2[4]), .c(n1467), .d(N314), 
        .out(n56) );
  inv U60 ( .in(n57), .out(n1083) );
  aoi22 U61 ( .a(n1505), .b(final_floor_elevator2[49]), .c(n1466), .d(N359), 
        .out(n57) );
  inv U62 ( .in(n58), .out(n1082) );
  aoi22 U63 ( .a(n1505), .b(final_floor_elevator2[48]), .c(n1466), .d(N358), 
        .out(n58) );
  inv U64 ( .in(n59), .out(n1081) );
  aoi22 U65 ( .a(n1505), .b(final_floor_elevator2[47]), .c(n1466), .d(N357), 
        .out(n59) );
  inv U66 ( .in(n60), .out(n1080) );
  aoi22 U67 ( .a(n1505), .b(final_floor_elevator2[46]), .c(n1465), .d(N356), 
        .out(n60) );
  inv U68 ( .in(n61), .out(n1079) );
  aoi22 U69 ( .a(n1505), .b(final_floor_elevator2[45]), .c(n1465), .d(N355), 
        .out(n61) );
  inv U70 ( .in(n62), .out(n1078) );
  aoi22 U71 ( .a(n1505), .b(final_floor_elevator2[44]), .c(n1465), .d(N354), 
        .out(n62) );
  inv U72 ( .in(n63), .out(n1077) );
  aoi22 U73 ( .a(n1505), .b(final_floor_elevator2[43]), .c(n1464), .d(N353), 
        .out(n63) );
  inv U74 ( .in(n64), .out(n1076) );
  aoi22 U75 ( .a(n1505), .b(final_floor_elevator2[42]), .c(n1464), .d(N352), 
        .out(n64) );
  inv U76 ( .in(n65), .out(n1075) );
  aoi22 U77 ( .a(n1504), .b(final_floor_elevator2[41]), .c(n1464), .d(N351), 
        .out(n65) );
  inv U78 ( .in(n66), .out(n1074) );
  aoi22 U79 ( .a(n1504), .b(final_floor_elevator2[40]), .c(n1463), .d(N350), 
        .out(n66) );
  inv U80 ( .in(n67), .out(n1037) );
  aoi22 U81 ( .a(n1504), .b(final_floor_elevator2[3]), .c(n1463), .d(N313), 
        .out(n67) );
  inv U82 ( .in(n68), .out(n1073) );
  aoi22 U83 ( .a(n1504), .b(final_floor_elevator2[39]), .c(n1463), .d(N349), 
        .out(n68) );
  inv U84 ( .in(n69), .out(n1072) );
  aoi22 U85 ( .a(n1504), .b(final_floor_elevator2[38]), .c(n1462), .d(N348), 
        .out(n69) );
  inv U86 ( .in(n70), .out(n1071) );
  aoi22 U87 ( .a(n1504), .b(final_floor_elevator2[37]), .c(n1462), .d(N347), 
        .out(n70) );
  inv U88 ( .in(n71), .out(n1070) );
  aoi22 U89 ( .a(n1504), .b(final_floor_elevator2[36]), .c(n1462), .d(N346), 
        .out(n71) );
  inv U90 ( .in(n72), .out(n1069) );
  aoi22 U91 ( .a(n1504), .b(final_floor_elevator2[35]), .c(n1461), .d(N345), 
        .out(n72) );
  inv U92 ( .in(n73), .out(n1068) );
  aoi22 U93 ( .a(n1504), .b(final_floor_elevator2[34]), .c(n1461), .d(N344), 
        .out(n73) );
  inv U94 ( .in(n74), .out(n1067) );
  aoi22 U95 ( .a(n1504), .b(final_floor_elevator2[33]), .c(n1461), .d(N343), 
        .out(n74) );
  inv U96 ( .in(n75), .out(n1066) );
  aoi22 U97 ( .a(n1504), .b(final_floor_elevator2[32]), .c(n1460), .d(N342), 
        .out(n75) );
  inv U98 ( .in(n76), .out(n1065) );
  aoi22 U99 ( .a(n1504), .b(final_floor_elevator2[31]), .c(n1460), .d(N341), 
        .out(n76) );
  inv U100 ( .in(n77), .out(n1064) );
  aoi22 U101 ( .a(n1503), .b(final_floor_elevator2[30]), .c(n1460), .d(N340), 
        .out(n77) );
  inv U102 ( .in(n78), .out(n1036) );
  aoi22 U103 ( .a(n1503), .b(final_floor_elevator2[2]), .c(n1459), .d(N312), 
        .out(n78) );
  inv U104 ( .in(n79), .out(n1063) );
  aoi22 U105 ( .a(n1503), .b(final_floor_elevator2[29]), .c(n1459), .d(N339), 
        .out(n79) );
  inv U106 ( .in(n80), .out(n1062) );
  aoi22 U107 ( .a(n1503), .b(final_floor_elevator2[28]), .c(n1459), .d(N338), 
        .out(n80) );
  inv U108 ( .in(n81), .out(n1061) );
  aoi22 U109 ( .a(n1503), .b(final_floor_elevator2[27]), .c(n1458), .d(N337), 
        .out(n81) );
  inv U110 ( .in(n82), .out(n1060) );
  aoi22 U111 ( .a(n1503), .b(final_floor_elevator2[26]), .c(n1458), .d(N336), 
        .out(n82) );
  inv U112 ( .in(n83), .out(n1059) );
  aoi22 U113 ( .a(n1503), .b(final_floor_elevator2[25]), .c(n1458), .d(N335), 
        .out(n83) );
  inv U114 ( .in(n84), .out(n1058) );
  aoi22 U115 ( .a(n1503), .b(final_floor_elevator2[24]), .c(n1457), .d(N334), 
        .out(n84) );
  inv U116 ( .in(n85), .out(n1057) );
  aoi22 U117 ( .a(n1503), .b(final_floor_elevator2[23]), .c(n1457), .d(N333), 
        .out(n85) );
  inv U118 ( .in(n86), .out(n1056) );
  aoi22 U119 ( .a(n1503), .b(final_floor_elevator2[22]), .c(n1457), .d(N332), 
        .out(n86) );
  inv U120 ( .in(n87), .out(n1055) );
  aoi22 U121 ( .a(n1503), .b(final_floor_elevator2[21]), .c(n1456), .d(N331), 
        .out(n87) );
  inv U122 ( .in(n88), .out(n1054) );
  aoi22 U123 ( .a(n1503), .b(final_floor_elevator2[20]), .c(n1456), .d(N330), 
        .out(n88) );
  inv U124 ( .in(n89), .out(n1035) );
  aoi22 U125 ( .a(n1502), .b(final_floor_elevator2[1]), .c(n1456), .d(N311), 
        .out(n89) );
  inv U126 ( .in(n90), .out(n1053) );
  aoi22 U127 ( .a(n1502), .b(final_floor_elevator2[19]), .c(n1455), .d(N329), 
        .out(n90) );
  inv U128 ( .in(n91), .out(n1052) );
  aoi22 U129 ( .a(n1502), .b(final_floor_elevator2[18]), .c(n1455), .d(N328), 
        .out(n91) );
  inv U130 ( .in(n92), .out(n1051) );
  aoi22 U131 ( .a(n1502), .b(final_floor_elevator2[17]), .c(n1455), .d(N327), 
        .out(n92) );
  inv U132 ( .in(n93), .out(n1050) );
  aoi22 U133 ( .a(n1502), .b(final_floor_elevator2[16]), .c(n1454), .d(N326), 
        .out(n93) );
  inv U134 ( .in(n94), .out(n1049) );
  aoi22 U135 ( .a(n1502), .b(final_floor_elevator2[15]), .c(n1454), .d(N325), 
        .out(n94) );
  inv U136 ( .in(n95), .out(n1048) );
  aoi22 U137 ( .a(n1502), .b(final_floor_elevator2[14]), .c(n1454), .d(N324), 
        .out(n95) );
  inv U138 ( .in(n96), .out(n1047) );
  aoi22 U139 ( .a(n1502), .b(final_floor_elevator2[13]), .c(n1453), .d(N323), 
        .out(n96) );
  inv U140 ( .in(n97), .out(n1046) );
  aoi22 U141 ( .a(n1502), .b(final_floor_elevator2[12]), .c(n1453), .d(N322), 
        .out(n97) );
  inv U142 ( .in(n98), .out(n1045) );
  aoi22 U143 ( .a(n1502), .b(final_floor_elevator2[11]), .c(n1453), .d(N321), 
        .out(n98) );
  inv U144 ( .in(n99), .out(n1044) );
  aoi22 U145 ( .a(n1502), .b(final_floor_elevator2[10]), .c(n1452), .d(N320), 
        .out(n99) );
  inv U146 ( .in(n100), .out(n1034) );
  aoi22 U147 ( .a(n1502), .b(final_floor_elevator2[0]), .c(n1452), .d(N310), 
        .out(n100) );
  inv U149 ( .in(n101), .out(n1107) );
  aoi22 U150 ( .a(n1589), .b(final_floor_elevator1[9]), .c(n1555), .d(N35), 
        .out(n101) );
  inv U151 ( .in(n102), .out(n1106) );
  aoi22 U152 ( .a(n1589), .b(final_floor_elevator1[8]), .c(n1555), .d(N34), 
        .out(n102) );
  inv U153 ( .in(n103), .out(n1105) );
  aoi22 U154 ( .a(n1589), .b(final_floor_elevator1[7]), .c(n1554), .d(N33), 
        .out(n103) );
  inv U155 ( .in(n104), .out(n1104) );
  aoi22 U156 ( .a(n1589), .b(final_floor_elevator1[6]), .c(n1554), .d(N32), 
        .out(n104) );
  inv U157 ( .in(n105), .out(n1148) );
  aoi22 U158 ( .a(n1554), .b(N90), .c(n1588), .d(\ne_47/SA ), .out(n105) );
  inv U159 ( .in(n106), .out(n1149) );
  aoi22 U160 ( .a(n1553), .b(N89), .c(n1588), .d(final_floor_elevator1[62]), 
        .out(n106) );
  inv U161 ( .in(n107), .out(n1150) );
  aoi22 U162 ( .a(n1553), .b(N88), .c(n1588), .d(final_floor_elevator1[61]), 
        .out(n107) );
  inv U163 ( .in(n108), .out(n1151) );
  aoi22 U164 ( .a(n1553), .b(N87), .c(n1588), .d(final_floor_elevator1[60]), 
        .out(n108) );
  inv U165 ( .in(n109), .out(n1103) );
  aoi22 U166 ( .a(n1588), .b(final_floor_elevator1[5]), .c(n1552), .d(N31), 
        .out(n109) );
  inv U167 ( .in(n110), .out(n1152) );
  aoi22 U168 ( .a(n1552), .b(N86), .c(n1588), .d(final_floor_elevator1[59]), 
        .out(n110) );
  inv U169 ( .in(n111), .out(n1153) );
  aoi22 U170 ( .a(n1552), .b(N85), .c(n1588), .d(final_floor_elevator1[58]), 
        .out(n111) );
  inv U171 ( .in(n112), .out(n1154) );
  aoi22 U172 ( .a(n1551), .b(N84), .c(n1588), .d(final_floor_elevator1[57]), 
        .out(n112) );
  inv U173 ( .in(n113), .out(n1155) );
  aoi22 U174 ( .a(n1551), .b(N83), .c(n1588), .d(final_floor_elevator1[56]), 
        .out(n113) );
  inv U175 ( .in(n114), .out(n1156) );
  aoi22 U176 ( .a(n1551), .b(N82), .c(n1588), .d(final_floor_elevator1[55]), 
        .out(n114) );
  inv U177 ( .in(n115), .out(n1157) );
  aoi22 U178 ( .a(n1550), .b(N81), .c(n1588), .d(final_floor_elevator1[54]), 
        .out(n115) );
  inv U179 ( .in(n116), .out(n1158) );
  aoi22 U180 ( .a(n1550), .b(N80), .c(n1588), .d(final_floor_elevator1[53]), 
        .out(n116) );
  inv U181 ( .in(n117), .out(n1159) );
  aoi22 U182 ( .a(n1550), .b(N79), .c(n1587), .d(final_floor_elevator1[52]), 
        .out(n117) );
  inv U183 ( .in(n118), .out(n1160) );
  aoi22 U184 ( .a(n1549), .b(N78), .c(n1587), .d(final_floor_elevator1[51]), 
        .out(n118) );
  inv U185 ( .in(n119), .out(n1161) );
  aoi22 U186 ( .a(n1549), .b(N77), .c(n1587), .d(final_floor_elevator1[50]), 
        .out(n119) );
  inv U187 ( .in(n120), .out(n1102) );
  aoi22 U188 ( .a(n1587), .b(final_floor_elevator1[4]), .c(n1549), .d(N30), 
        .out(n120) );
  inv U189 ( .in(n121), .out(n1147) );
  aoi22 U190 ( .a(n1587), .b(final_floor_elevator1[49]), .c(n1548), .d(N75), 
        .out(n121) );
  inv U191 ( .in(n122), .out(n1146) );
  aoi22 U192 ( .a(n1587), .b(final_floor_elevator1[48]), .c(n1548), .d(N74), 
        .out(n122) );
  inv U193 ( .in(n123), .out(n1145) );
  aoi22 U194 ( .a(n1587), .b(final_floor_elevator1[47]), .c(n1548), .d(N73), 
        .out(n123) );
  inv U195 ( .in(n124), .out(n1144) );
  aoi22 U196 ( .a(n1587), .b(final_floor_elevator1[46]), .c(n1547), .d(N72), 
        .out(n124) );
  inv U197 ( .in(n125), .out(n1143) );
  aoi22 U198 ( .a(n1587), .b(final_floor_elevator1[45]), .c(n1547), .d(N71), 
        .out(n125) );
  inv U199 ( .in(n126), .out(n1142) );
  aoi22 U200 ( .a(n1587), .b(final_floor_elevator1[44]), .c(n1547), .d(N70), 
        .out(n126) );
  inv U201 ( .in(n127), .out(n1141) );
  aoi22 U202 ( .a(n1587), .b(final_floor_elevator1[43]), .c(n1546), .d(N69), 
        .out(n127) );
  inv U203 ( .in(n128), .out(n1140) );
  aoi22 U204 ( .a(n1587), .b(final_floor_elevator1[42]), .c(n1546), .d(N68), 
        .out(n128) );
  inv U205 ( .in(n129), .out(n1139) );
  aoi22 U206 ( .a(n1586), .b(final_floor_elevator1[41]), .c(n1546), .d(N67), 
        .out(n129) );
  inv U207 ( .in(n130), .out(n1138) );
  aoi22 U208 ( .a(n1586), .b(final_floor_elevator1[40]), .c(n1545), .d(N66), 
        .out(n130) );
  inv U209 ( .in(n131), .out(n1101) );
  aoi22 U210 ( .a(n1586), .b(final_floor_elevator1[3]), .c(n1545), .d(N29), 
        .out(n131) );
  inv U211 ( .in(n132), .out(n1137) );
  aoi22 U212 ( .a(n1586), .b(final_floor_elevator1[39]), .c(n1545), .d(N65), 
        .out(n132) );
  inv U213 ( .in(n133), .out(n1136) );
  aoi22 U214 ( .a(n1586), .b(final_floor_elevator1[38]), .c(n1544), .d(N64), 
        .out(n133) );
  inv U215 ( .in(n134), .out(n1135) );
  aoi22 U216 ( .a(n1586), .b(final_floor_elevator1[37]), .c(n1544), .d(N63), 
        .out(n134) );
  inv U217 ( .in(n135), .out(n1134) );
  aoi22 U218 ( .a(n1586), .b(final_floor_elevator1[36]), .c(n1544), .d(N62), 
        .out(n135) );
  inv U219 ( .in(n136), .out(n1133) );
  aoi22 U220 ( .a(n1586), .b(final_floor_elevator1[35]), .c(n1543), .d(N61), 
        .out(n136) );
  inv U221 ( .in(n137), .out(n1132) );
  aoi22 U222 ( .a(n1586), .b(final_floor_elevator1[34]), .c(n1543), .d(N60), 
        .out(n137) );
  inv U223 ( .in(n138), .out(n1131) );
  aoi22 U224 ( .a(n1586), .b(final_floor_elevator1[33]), .c(n1543), .d(N59), 
        .out(n138) );
  inv U225 ( .in(n139), .out(n1130) );
  aoi22 U226 ( .a(n1586), .b(final_floor_elevator1[32]), .c(n1542), .d(N58), 
        .out(n139) );
  inv U227 ( .in(n140), .out(n1129) );
  aoi22 U228 ( .a(n1586), .b(final_floor_elevator1[31]), .c(n1542), .d(N57), 
        .out(n140) );
  inv U229 ( .in(n141), .out(n1128) );
  aoi22 U230 ( .a(n1585), .b(final_floor_elevator1[30]), .c(n1542), .d(N56), 
        .out(n141) );
  inv U231 ( .in(n142), .out(n1100) );
  aoi22 U232 ( .a(n1585), .b(final_floor_elevator1[2]), .c(n1541), .d(N28), 
        .out(n142) );
  inv U233 ( .in(n143), .out(n1127) );
  aoi22 U234 ( .a(n1585), .b(final_floor_elevator1[29]), .c(n1541), .d(N55), 
        .out(n143) );
  inv U235 ( .in(n144), .out(n1126) );
  aoi22 U236 ( .a(n1585), .b(final_floor_elevator1[28]), .c(n1541), .d(N54), 
        .out(n144) );
  inv U237 ( .in(n145), .out(n1125) );
  aoi22 U238 ( .a(n1585), .b(final_floor_elevator1[27]), .c(n1540), .d(N53), 
        .out(n145) );
  inv U239 ( .in(n146), .out(n1124) );
  aoi22 U240 ( .a(n1585), .b(final_floor_elevator1[26]), .c(n1540), .d(N52), 
        .out(n146) );
  inv U241 ( .in(n147), .out(n1123) );
  aoi22 U242 ( .a(n1585), .b(final_floor_elevator1[25]), .c(n1540), .d(N51), 
        .out(n147) );
  inv U243 ( .in(n148), .out(n1122) );
  aoi22 U244 ( .a(n1585), .b(final_floor_elevator1[24]), .c(n1539), .d(N50), 
        .out(n148) );
  inv U245 ( .in(n149), .out(n1121) );
  aoi22 U246 ( .a(n1585), .b(final_floor_elevator1[23]), .c(n1539), .d(N49), 
        .out(n149) );
  inv U247 ( .in(n150), .out(n1120) );
  aoi22 U248 ( .a(n1585), .b(final_floor_elevator1[22]), .c(n1539), .d(N48), 
        .out(n150) );
  inv U249 ( .in(n151), .out(n1119) );
  aoi22 U250 ( .a(n1585), .b(final_floor_elevator1[21]), .c(n1538), .d(N47), 
        .out(n151) );
  inv U251 ( .in(n152), .out(n1118) );
  aoi22 U252 ( .a(n1585), .b(final_floor_elevator1[20]), .c(n1538), .d(N46), 
        .out(n152) );
  inv U253 ( .in(n153), .out(n1099) );
  aoi22 U254 ( .a(n1584), .b(final_floor_elevator1[1]), .c(n1538), .d(N27), 
        .out(n153) );
  inv U255 ( .in(n154), .out(n1117) );
  aoi22 U256 ( .a(n1584), .b(final_floor_elevator1[19]), .c(n1537), .d(N45), 
        .out(n154) );
  inv U257 ( .in(n155), .out(n1116) );
  aoi22 U258 ( .a(n1584), .b(final_floor_elevator1[18]), .c(n1537), .d(N44), 
        .out(n155) );
  inv U259 ( .in(n156), .out(n1115) );
  aoi22 U260 ( .a(n1584), .b(final_floor_elevator1[17]), .c(n1537), .d(N43), 
        .out(n156) );
  inv U261 ( .in(n157), .out(n1114) );
  aoi22 U262 ( .a(n1584), .b(final_floor_elevator1[16]), .c(n1536), .d(N42), 
        .out(n157) );
  inv U263 ( .in(n158), .out(n1113) );
  aoi22 U264 ( .a(n1584), .b(final_floor_elevator1[15]), .c(n1536), .d(N41), 
        .out(n158) );
  inv U265 ( .in(n159), .out(n1112) );
  aoi22 U266 ( .a(n1584), .b(final_floor_elevator1[14]), .c(n1536), .d(N40), 
        .out(n159) );
  inv U267 ( .in(n160), .out(n1111) );
  aoi22 U268 ( .a(n1584), .b(final_floor_elevator1[13]), .c(n1535), .d(N39), 
        .out(n160) );
  inv U269 ( .in(n161), .out(n1110) );
  aoi22 U270 ( .a(n1584), .b(final_floor_elevator1[12]), .c(n1535), .d(N38), 
        .out(n161) );
  inv U271 ( .in(n162), .out(n1109) );
  aoi22 U272 ( .a(n1584), .b(final_floor_elevator1[11]), .c(n1535), .d(N37), 
        .out(n162) );
  inv U273 ( .in(n163), .out(n1108) );
  aoi22 U274 ( .a(n1584), .b(final_floor_elevator1[10]), .c(n1534), .d(N36), 
        .out(n163) );
  inv U275 ( .in(n164), .out(n1098) );
  aoi22 U276 ( .a(n1584), .b(final_floor_elevator1[0]), .c(n1534), .d(N26), 
        .out(n164) );
  nand3 U278 ( .a(n26), .b(n1168), .c(n165), .out(n969) );
  nand3 U279 ( .a(n32), .b(n1618), .c(elevator2_status), .out(n165) );
  nand3 U280 ( .a(n23), .b(n1166), .c(n166), .out(n901) );
  nand3 U281 ( .a(n167), .b(n1663), .c(elevator1_status), .out(n166) );
  nand2 U282 ( .a(n26), .b(n169), .out(n968) );
  nand3 U283 ( .a(n170), .b(n1168), .c(direction_elevator2[1]), .out(n169) );
  nand2 U284 ( .a(n1168), .b(n171), .out(n966) );
  nand3 U285 ( .a(n170), .b(n26), .c(direction_elevator2[0]), .out(n171) );
  inv U286 ( .in(n172), .out(n26) );
  nor3 U287 ( .a(in_emergency_elevator2), .b(n1595), .c(n173), .out(n170) );
  inv U288 ( .in(n32), .out(n173) );
  nand2 U289 ( .a(n23), .b(n174), .out(n900) );
  nand3 U290 ( .a(n175), .b(n1166), .c(direction_elevator1[1]), .out(n174) );
  nand2 U291 ( .a(n1166), .b(n176), .out(n898) );
  nand3 U292 ( .a(n175), .b(n23), .c(direction_elevator1[0]), .out(n176) );
  inv U293 ( .in(n177), .out(n23) );
  nor3 U294 ( .a(in_emergency_elevator1), .b(n1640), .c(n35), .out(n175) );
  inv U295 ( .in(n167), .out(n35) );
  nand2 U296 ( .a(n178), .b(n179), .out(n1024) );
  aoi22 U297 ( .a(n172), .b(N428), .c(N430), .d(n180), .out(n179) );
  aoi22 U298 ( .a(current_floor_elevator2[9]), .b(n181), .c(
        current_floor_output_elevator2[9]), .d(n182), .out(n178) );
  nand2 U299 ( .a(n183), .b(n184), .out(n1025) );
  aoi22 U300 ( .a(n172), .b(N429), .c(N431), .d(n180), .out(n184) );
  aoi22 U301 ( .a(current_floor_elevator2[8]), .b(n181), .c(
        current_floor_output_elevator2[8]), .d(n182), .out(n183) );
  nand2 U302 ( .a(n185), .b(n186), .out(n1026) );
  aoi22 U303 ( .a(n172), .b(N430), .c(N432), .d(n180), .out(n186) );
  aoi22 U304 ( .a(current_floor_elevator2[7]), .b(n181), .c(
        current_floor_output_elevator2[7]), .d(n182), .out(n185) );
  nand2 U305 ( .a(n187), .b(n188), .out(n1027) );
  aoi22 U306 ( .a(n172), .b(N431), .c(N433), .d(n180), .out(n188) );
  aoi22 U307 ( .a(current_floor_elevator2[6]), .b(n181), .c(
        current_floor_output_elevator2[6]), .d(n182), .out(n187) );
  nand2 U308 ( .a(n189), .b(n190), .out(n970) );
  nand2 U309 ( .a(\eq_47_3/SA ), .b(n182), .out(n190) );
  aoi22 U310 ( .a(N376), .b(n180), .c(current_floor_elevator2[63]), .d(n181), 
        .out(n189) );
  nand2 U311 ( .a(n191), .b(n192), .out(n971) );
  aoi22 U312 ( .a(n172), .b(\r126/SB ), .c(N377), .d(n180), .out(n192) );
  aoi22 U313 ( .a(current_floor_elevator2[62]), .b(n181), .c(
        current_floor_output_elevator2[62]), .d(n182), .out(n191) );
  nand2 U314 ( .a(n193), .b(n194), .out(n972) );
  aoi22 U315 ( .a(n172), .b(N376), .c(N378), .d(n180), .out(n194) );
  aoi22 U316 ( .a(current_floor_elevator2[61]), .b(n181), .c(
        current_floor_output_elevator2[61]), .d(n182), .out(n193) );
  nand2 U317 ( .a(n195), .b(n196), .out(n973) );
  aoi22 U318 ( .a(n172), .b(N377), .c(N379), .d(n180), .out(n196) );
  aoi22 U319 ( .a(current_floor_elevator2[60]), .b(n181), .c(
        current_floor_output_elevator2[60]), .d(n182), .out(n195) );
  nand2 U320 ( .a(n197), .b(n198), .out(n1028) );
  aoi22 U321 ( .a(n172), .b(N432), .c(N434), .d(n180), .out(n198) );
  aoi22 U322 ( .a(current_floor_elevator2[5]), .b(n181), .c(
        current_floor_output_elevator2[5]), .d(n182), .out(n197) );
  nand2 U323 ( .a(n199), .b(n200), .out(n974) );
  aoi22 U324 ( .a(n172), .b(N378), .c(N380), .d(n180), .out(n200) );
  aoi22 U325 ( .a(current_floor_elevator2[59]), .b(n181), .c(
        current_floor_output_elevator2[59]), .d(n182), .out(n199) );
  nand2 U326 ( .a(n201), .b(n202), .out(n975) );
  aoi22 U327 ( .a(n172), .b(N379), .c(N381), .d(n180), .out(n202) );
  aoi22 U328 ( .a(current_floor_elevator2[58]), .b(n181), .c(
        current_floor_output_elevator2[58]), .d(n182), .out(n201) );
  nand2 U329 ( .a(n203), .b(n204), .out(n976) );
  aoi22 U330 ( .a(n172), .b(N380), .c(N382), .d(n180), .out(n204) );
  aoi22 U331 ( .a(current_floor_elevator2[57]), .b(n181), .c(
        current_floor_output_elevator2[57]), .d(n182), .out(n203) );
  nand2 U332 ( .a(n205), .b(n206), .out(n977) );
  aoi22 U333 ( .a(n172), .b(N381), .c(N383), .d(n180), .out(n206) );
  aoi22 U334 ( .a(current_floor_elevator2[56]), .b(n181), .c(
        current_floor_output_elevator2[56]), .d(n182), .out(n205) );
  nand2 U335 ( .a(n207), .b(n208), .out(n978) );
  aoi22 U336 ( .a(n172), .b(N382), .c(N384), .d(n180), .out(n208) );
  aoi22 U337 ( .a(current_floor_elevator2[55]), .b(n181), .c(
        current_floor_output_elevator2[55]), .d(n182), .out(n207) );
  nand2 U338 ( .a(n209), .b(n210), .out(n979) );
  aoi22 U339 ( .a(n172), .b(N383), .c(N385), .d(n180), .out(n210) );
  aoi22 U340 ( .a(current_floor_elevator2[54]), .b(n181), .c(
        current_floor_output_elevator2[54]), .d(n182), .out(n209) );
  nand2 U341 ( .a(n211), .b(n212), .out(n980) );
  aoi22 U342 ( .a(n172), .b(N384), .c(N386), .d(n180), .out(n212) );
  aoi22 U343 ( .a(current_floor_elevator2[53]), .b(n181), .c(
        current_floor_output_elevator2[53]), .d(n182), .out(n211) );
  nand2 U344 ( .a(n213), .b(n214), .out(n981) );
  aoi22 U345 ( .a(n172), .b(N385), .c(N387), .d(n180), .out(n214) );
  aoi22 U346 ( .a(current_floor_elevator2[52]), .b(n181), .c(
        current_floor_output_elevator2[52]), .d(n182), .out(n213) );
  nand2 U347 ( .a(n215), .b(n216), .out(n982) );
  aoi22 U348 ( .a(n172), .b(N386), .c(N388), .d(n180), .out(n216) );
  aoi22 U349 ( .a(current_floor_elevator2[51]), .b(n181), .c(
        current_floor_output_elevator2[51]), .d(n182), .out(n215) );
  nand2 U350 ( .a(n217), .b(n218), .out(n983) );
  aoi22 U351 ( .a(n172), .b(N387), .c(N389), .d(n180), .out(n218) );
  aoi22 U352 ( .a(current_floor_elevator2[50]), .b(n181), .c(
        current_floor_output_elevator2[50]), .d(n182), .out(n217) );
  nand2 U353 ( .a(n219), .b(n220), .out(n1029) );
  aoi22 U354 ( .a(n172), .b(N433), .c(N435), .d(n180), .out(n220) );
  aoi22 U355 ( .a(current_floor_elevator2[4]), .b(n181), .c(
        current_floor_output_elevator2[4]), .d(n182), .out(n219) );
  nand2 U356 ( .a(n221), .b(n222), .out(n984) );
  aoi22 U357 ( .a(n172), .b(N388), .c(N390), .d(n180), .out(n222) );
  aoi22 U358 ( .a(current_floor_elevator2[49]), .b(n181), .c(
        current_floor_output_elevator2[49]), .d(n182), .out(n221) );
  nand2 U359 ( .a(n223), .b(n224), .out(n985) );
  aoi22 U360 ( .a(n172), .b(N389), .c(N391), .d(n180), .out(n224) );
  aoi22 U361 ( .a(current_floor_elevator2[48]), .b(n181), .c(
        current_floor_output_elevator2[48]), .d(n182), .out(n223) );
  nand2 U362 ( .a(n225), .b(n226), .out(n986) );
  aoi22 U363 ( .a(n172), .b(N390), .c(N392), .d(n180), .out(n226) );
  aoi22 U364 ( .a(current_floor_elevator2[47]), .b(n181), .c(
        current_floor_output_elevator2[47]), .d(n182), .out(n225) );
  nand2 U365 ( .a(n227), .b(n228), .out(n987) );
  aoi22 U366 ( .a(n172), .b(N391), .c(N393), .d(n180), .out(n228) );
  aoi22 U367 ( .a(current_floor_elevator2[46]), .b(n181), .c(
        current_floor_output_elevator2[46]), .d(n182), .out(n227) );
  nand2 U368 ( .a(n229), .b(n230), .out(n988) );
  aoi22 U369 ( .a(n172), .b(N392), .c(N394), .d(n180), .out(n230) );
  aoi22 U370 ( .a(current_floor_elevator2[45]), .b(n181), .c(
        current_floor_output_elevator2[45]), .d(n182), .out(n229) );
  nand2 U371 ( .a(n231), .b(n232), .out(n989) );
  aoi22 U372 ( .a(n172), .b(N393), .c(N395), .d(n180), .out(n232) );
  aoi22 U373 ( .a(current_floor_elevator2[44]), .b(n181), .c(
        current_floor_output_elevator2[44]), .d(n182), .out(n231) );
  nand2 U374 ( .a(n233), .b(n234), .out(n990) );
  aoi22 U375 ( .a(n172), .b(N394), .c(N396), .d(n180), .out(n234) );
  aoi22 U376 ( .a(current_floor_elevator2[43]), .b(n181), .c(
        current_floor_output_elevator2[43]), .d(n182), .out(n233) );
  nand2 U377 ( .a(n235), .b(n236), .out(n991) );
  aoi22 U378 ( .a(n172), .b(N395), .c(N397), .d(n180), .out(n236) );
  aoi22 U379 ( .a(current_floor_elevator2[42]), .b(n181), .c(
        current_floor_output_elevator2[42]), .d(n182), .out(n235) );
  nand2 U380 ( .a(n237), .b(n238), .out(n992) );
  aoi22 U381 ( .a(n172), .b(N396), .c(N398), .d(n180), .out(n238) );
  aoi22 U382 ( .a(current_floor_elevator2[41]), .b(n181), .c(
        current_floor_output_elevator2[41]), .d(n182), .out(n237) );
  nand2 U383 ( .a(n239), .b(n240), .out(n993) );
  aoi22 U384 ( .a(n172), .b(N397), .c(N399), .d(n180), .out(n240) );
  aoi22 U385 ( .a(current_floor_elevator2[40]), .b(n181), .c(
        current_floor_output_elevator2[40]), .d(n182), .out(n239) );
  nand2 U386 ( .a(n241), .b(n242), .out(n1030) );
  aoi22 U387 ( .a(n172), .b(N434), .c(N436), .d(n180), .out(n242) );
  aoi22 U388 ( .a(current_floor_elevator2[3]), .b(n181), .c(
        current_floor_output_elevator2[3]), .d(n182), .out(n241) );
  nand2 U389 ( .a(n243), .b(n244), .out(n994) );
  aoi22 U390 ( .a(n172), .b(N398), .c(N400), .d(n180), .out(n244) );
  aoi22 U391 ( .a(current_floor_elevator2[39]), .b(n181), .c(
        current_floor_output_elevator2[39]), .d(n182), .out(n243) );
  nand2 U392 ( .a(n245), .b(n246), .out(n995) );
  aoi22 U393 ( .a(n172), .b(N399), .c(N401), .d(n180), .out(n246) );
  aoi22 U394 ( .a(current_floor_elevator2[38]), .b(n181), .c(
        current_floor_output_elevator2[38]), .d(n182), .out(n245) );
  nand2 U395 ( .a(n247), .b(n248), .out(n996) );
  aoi22 U396 ( .a(n172), .b(N400), .c(N402), .d(n180), .out(n248) );
  aoi22 U397 ( .a(current_floor_elevator2[37]), .b(n181), .c(
        current_floor_output_elevator2[37]), .d(n182), .out(n247) );
  nand2 U398 ( .a(n249), .b(n250), .out(n997) );
  aoi22 U399 ( .a(n172), .b(N401), .c(N403), .d(n180), .out(n250) );
  aoi22 U400 ( .a(current_floor_elevator2[36]), .b(n181), .c(
        current_floor_output_elevator2[36]), .d(n182), .out(n249) );
  nand2 U401 ( .a(n251), .b(n252), .out(n998) );
  aoi22 U402 ( .a(n172), .b(N402), .c(N404), .d(n180), .out(n252) );
  aoi22 U403 ( .a(current_floor_elevator2[35]), .b(n181), .c(
        current_floor_output_elevator2[35]), .d(n182), .out(n251) );
  nand2 U404 ( .a(n253), .b(n254), .out(n999) );
  aoi22 U405 ( .a(n172), .b(N403), .c(N405), .d(n180), .out(n254) );
  aoi22 U406 ( .a(current_floor_elevator2[34]), .b(n181), .c(
        current_floor_output_elevator2[34]), .d(n182), .out(n253) );
  nand2 U407 ( .a(n255), .b(n256), .out(n1000) );
  aoi22 U408 ( .a(n172), .b(N404), .c(N406), .d(n180), .out(n256) );
  aoi22 U409 ( .a(current_floor_elevator2[33]), .b(n181), .c(
        current_floor_output_elevator2[33]), .d(n182), .out(n255) );
  nand2 U410 ( .a(n257), .b(n258), .out(n1001) );
  aoi22 U411 ( .a(n172), .b(N405), .c(N407), .d(n180), .out(n258) );
  aoi22 U412 ( .a(current_floor_elevator2[32]), .b(n181), .c(
        current_floor_output_elevator2[32]), .d(n182), .out(n257) );
  nand2 U413 ( .a(n259), .b(n260), .out(n1002) );
  aoi22 U414 ( .a(n172), .b(N406), .c(N408), .d(n180), .out(n260) );
  aoi22 U415 ( .a(current_floor_elevator2[31]), .b(n181), .c(
        current_floor_output_elevator2[31]), .d(n182), .out(n259) );
  nand2 U416 ( .a(n261), .b(n262), .out(n1003) );
  aoi22 U417 ( .a(n172), .b(N407), .c(N409), .d(n180), .out(n262) );
  aoi22 U418 ( .a(current_floor_elevator2[30]), .b(n181), .c(
        current_floor_output_elevator2[30]), .d(n182), .out(n261) );
  nand2 U419 ( .a(n263), .b(n264), .out(n1031) );
  aoi22 U420 ( .a(n172), .b(N435), .c(N437), .d(n180), .out(n264) );
  aoi22 U421 ( .a(current_floor_elevator2[2]), .b(n181), .c(
        current_floor_output_elevator2[2]), .d(n182), .out(n263) );
  nand2 U422 ( .a(n265), .b(n266), .out(n1004) );
  aoi22 U423 ( .a(n172), .b(N408), .c(N410), .d(n180), .out(n266) );
  aoi22 U424 ( .a(current_floor_elevator2[29]), .b(n181), .c(
        current_floor_output_elevator2[29]), .d(n182), .out(n265) );
  nand2 U425 ( .a(n267), .b(n268), .out(n1005) );
  aoi22 U426 ( .a(n172), .b(N409), .c(N411), .d(n180), .out(n268) );
  aoi22 U427 ( .a(current_floor_elevator2[28]), .b(n181), .c(
        current_floor_output_elevator2[28]), .d(n182), .out(n267) );
  nand2 U428 ( .a(n269), .b(n270), .out(n1006) );
  aoi22 U429 ( .a(n172), .b(N410), .c(N412), .d(n180), .out(n270) );
  aoi22 U430 ( .a(current_floor_elevator2[27]), .b(n181), .c(
        current_floor_output_elevator2[27]), .d(n182), .out(n269) );
  nand2 U431 ( .a(n271), .b(n272), .out(n1007) );
  aoi22 U432 ( .a(n172), .b(N411), .c(N413), .d(n180), .out(n272) );
  aoi22 U433 ( .a(current_floor_elevator2[26]), .b(n181), .c(
        current_floor_output_elevator2[26]), .d(n182), .out(n271) );
  nand2 U434 ( .a(n273), .b(n274), .out(n1008) );
  aoi22 U435 ( .a(n172), .b(N412), .c(N414), .d(n180), .out(n274) );
  aoi22 U436 ( .a(current_floor_elevator2[25]), .b(n181), .c(
        current_floor_output_elevator2[25]), .d(n182), .out(n273) );
  nand2 U437 ( .a(n275), .b(n276), .out(n1009) );
  aoi22 U438 ( .a(n172), .b(N413), .c(N415), .d(n180), .out(n276) );
  aoi22 U439 ( .a(current_floor_elevator2[24]), .b(n181), .c(
        current_floor_output_elevator2[24]), .d(n182), .out(n275) );
  nand2 U440 ( .a(n277), .b(n278), .out(n1010) );
  aoi22 U441 ( .a(n172), .b(N414), .c(N416), .d(n180), .out(n278) );
  aoi22 U442 ( .a(current_floor_elevator2[23]), .b(n181), .c(
        current_floor_output_elevator2[23]), .d(n182), .out(n277) );
  nand2 U443 ( .a(n279), .b(n280), .out(n1011) );
  aoi22 U444 ( .a(n172), .b(N415), .c(N417), .d(n180), .out(n280) );
  aoi22 U445 ( .a(current_floor_elevator2[22]), .b(n181), .c(
        current_floor_output_elevator2[22]), .d(n182), .out(n279) );
  nand2 U446 ( .a(n281), .b(n282), .out(n1012) );
  aoi22 U447 ( .a(n172), .b(N416), .c(N418), .d(n180), .out(n282) );
  aoi22 U448 ( .a(current_floor_elevator2[21]), .b(n181), .c(
        current_floor_output_elevator2[21]), .d(n182), .out(n281) );
  nand2 U449 ( .a(n283), .b(n284), .out(n1013) );
  aoi22 U450 ( .a(n172), .b(N417), .c(N419), .d(n180), .out(n284) );
  aoi22 U451 ( .a(current_floor_elevator2[20]), .b(n181), .c(
        current_floor_output_elevator2[20]), .d(n182), .out(n283) );
  nand2 U452 ( .a(n285), .b(n286), .out(n1032) );
  aoi22 U453 ( .a(n172), .b(N436), .c(N438), .d(n180), .out(n286) );
  aoi22 U454 ( .a(current_floor_elevator2[1]), .b(n181), .c(
        current_floor_output_elevator2[1]), .d(n182), .out(n285) );
  nand2 U455 ( .a(n287), .b(n288), .out(n1014) );
  aoi22 U456 ( .a(n172), .b(N418), .c(N420), .d(n180), .out(n288) );
  aoi22 U457 ( .a(current_floor_elevator2[19]), .b(n181), .c(
        current_floor_output_elevator2[19]), .d(n182), .out(n287) );
  nand2 U458 ( .a(n289), .b(n290), .out(n1015) );
  aoi22 U459 ( .a(n172), .b(N419), .c(N421), .d(n180), .out(n290) );
  aoi22 U460 ( .a(current_floor_elevator2[18]), .b(n181), .c(
        current_floor_output_elevator2[18]), .d(n182), .out(n289) );
  nand2 U461 ( .a(n291), .b(n292), .out(n1016) );
  aoi22 U462 ( .a(n172), .b(N420), .c(N422), .d(n180), .out(n292) );
  aoi22 U463 ( .a(current_floor_elevator2[17]), .b(n181), .c(
        current_floor_output_elevator2[17]), .d(n182), .out(n291) );
  nand2 U464 ( .a(n293), .b(n294), .out(n1017) );
  aoi22 U465 ( .a(n172), .b(N421), .c(N423), .d(n180), .out(n294) );
  aoi22 U466 ( .a(current_floor_elevator2[16]), .b(n181), .c(
        current_floor_output_elevator2[16]), .d(n182), .out(n293) );
  nand2 U467 ( .a(n295), .b(n296), .out(n1018) );
  aoi22 U468 ( .a(n172), .b(N422), .c(N424), .d(n180), .out(n296) );
  aoi22 U469 ( .a(current_floor_elevator2[15]), .b(n181), .c(
        current_floor_output_elevator2[15]), .d(n182), .out(n295) );
  nand2 U470 ( .a(n297), .b(n298), .out(n1019) );
  aoi22 U471 ( .a(n172), .b(N423), .c(N425), .d(n180), .out(n298) );
  aoi22 U472 ( .a(current_floor_elevator2[14]), .b(n181), .c(
        current_floor_output_elevator2[14]), .d(n182), .out(n297) );
  nand2 U473 ( .a(n299), .b(n300), .out(n1020) );
  aoi22 U474 ( .a(n172), .b(N424), .c(N426), .d(n180), .out(n300) );
  aoi22 U475 ( .a(current_floor_elevator2[13]), .b(n181), .c(
        current_floor_output_elevator2[13]), .d(n182), .out(n299) );
  nand2 U476 ( .a(n301), .b(n302), .out(n1021) );
  aoi22 U477 ( .a(n172), .b(N425), .c(N427), .d(n180), .out(n302) );
  aoi22 U478 ( .a(current_floor_elevator2[12]), .b(n181), .c(
        current_floor_output_elevator2[12]), .d(n182), .out(n301) );
  nand2 U479 ( .a(n303), .b(n304), .out(n1022) );
  aoi22 U480 ( .a(n172), .b(N426), .c(N428), .d(n180), .out(n304) );
  aoi22 U481 ( .a(current_floor_elevator2[11]), .b(n181), .c(
        current_floor_output_elevator2[11]), .d(n182), .out(n303) );
  nand2 U482 ( .a(n305), .b(n306), .out(n1023) );
  aoi22 U483 ( .a(n172), .b(N427), .c(N429), .d(n180), .out(n306) );
  aoi22 U484 ( .a(current_floor_elevator2[10]), .b(n181), .c(
        current_floor_output_elevator2[10]), .d(n182), .out(n305) );
  nand2 U485 ( .a(n307), .b(n308), .out(n1033) );
  nand2 U486 ( .a(current_floor_output_elevator2[0]), .b(n182), .out(n308) );
  aoi22 U487 ( .a(n172), .b(N437), .c(current_floor_elevator2[0]), .d(n181), 
        .out(n307) );
  nor2 U488 ( .a(n182), .b(n1170), .out(n181) );
  nand2 U489 ( .a(n309), .b(n310), .out(n956) );
  aoi22 U490 ( .a(n177), .b(N144), .c(N146), .d(n311), .out(n310) );
  aoi22 U491 ( .a(current_floor_elevator1[9]), .b(n312), .c(
        current_floor_output_elevator1[9]), .d(n313), .out(n309) );
  nand2 U492 ( .a(n314), .b(n315), .out(n957) );
  aoi22 U493 ( .a(n177), .b(N145), .c(N147), .d(n311), .out(n315) );
  aoi22 U494 ( .a(current_floor_elevator1[8]), .b(n312), .c(
        current_floor_output_elevator1[8]), .d(n313), .out(n314) );
  nand2 U495 ( .a(n316), .b(n317), .out(n958) );
  aoi22 U496 ( .a(n177), .b(N146), .c(N148), .d(n311), .out(n317) );
  aoi22 U497 ( .a(current_floor_elevator1[7]), .b(n312), .c(
        current_floor_output_elevator1[7]), .d(n313), .out(n316) );
  nand2 U498 ( .a(n318), .b(n319), .out(n959) );
  aoi22 U499 ( .a(n177), .b(N147), .c(N149), .d(n311), .out(n319) );
  aoi22 U500 ( .a(current_floor_elevator1[6]), .b(n312), .c(
        current_floor_output_elevator1[6]), .d(n313), .out(n318) );
  nand2 U501 ( .a(n320), .b(n321), .out(n902) );
  nand2 U502 ( .a(\eq_42_3/SA ), .b(n313), .out(n321) );
  aoi22 U503 ( .a(N92), .b(n311), .c(current_floor_elevator1[63]), .d(n312), 
        .out(n320) );
  nand2 U504 ( .a(n322), .b(n323), .out(n903) );
  aoi22 U505 ( .a(n177), .b(\r125/SB ), .c(N93), .d(n311), .out(n323) );
  aoi22 U506 ( .a(current_floor_elevator1[62]), .b(n312), .c(
        current_floor_output_elevator1[62]), .d(n313), .out(n322) );
  nand2 U507 ( .a(n324), .b(n325), .out(n904) );
  aoi22 U508 ( .a(n177), .b(N92), .c(N94), .d(n311), .out(n325) );
  aoi22 U509 ( .a(current_floor_elevator1[61]), .b(n312), .c(
        current_floor_output_elevator1[61]), .d(n313), .out(n324) );
  nand2 U510 ( .a(n326), .b(n327), .out(n905) );
  aoi22 U511 ( .a(n177), .b(N93), .c(N95), .d(n311), .out(n327) );
  aoi22 U512 ( .a(current_floor_elevator1[60]), .b(n312), .c(
        current_floor_output_elevator1[60]), .d(n313), .out(n326) );
  nand2 U513 ( .a(n328), .b(n329), .out(n960) );
  aoi22 U514 ( .a(n177), .b(N148), .c(N150), .d(n311), .out(n329) );
  aoi22 U515 ( .a(current_floor_elevator1[5]), .b(n312), .c(
        current_floor_output_elevator1[5]), .d(n313), .out(n328) );
  nand2 U516 ( .a(n330), .b(n331), .out(n906) );
  aoi22 U517 ( .a(n177), .b(N94), .c(N96), .d(n311), .out(n331) );
  aoi22 U518 ( .a(current_floor_elevator1[59]), .b(n312), .c(
        current_floor_output_elevator1[59]), .d(n313), .out(n330) );
  nand2 U519 ( .a(n332), .b(n333), .out(n907) );
  aoi22 U520 ( .a(n177), .b(N95), .c(N97), .d(n311), .out(n333) );
  aoi22 U521 ( .a(current_floor_elevator1[58]), .b(n312), .c(
        current_floor_output_elevator1[58]), .d(n313), .out(n332) );
  nand2 U522 ( .a(n334), .b(n335), .out(n908) );
  aoi22 U523 ( .a(n177), .b(N96), .c(N98), .d(n311), .out(n335) );
  aoi22 U524 ( .a(current_floor_elevator1[57]), .b(n312), .c(
        current_floor_output_elevator1[57]), .d(n313), .out(n334) );
  nand2 U525 ( .a(n336), .b(n337), .out(n909) );
  aoi22 U526 ( .a(n177), .b(N97), .c(N99), .d(n311), .out(n337) );
  aoi22 U527 ( .a(current_floor_elevator1[56]), .b(n312), .c(
        current_floor_output_elevator1[56]), .d(n313), .out(n336) );
  nand2 U528 ( .a(n338), .b(n339), .out(n910) );
  aoi22 U529 ( .a(n177), .b(N98), .c(N100), .d(n311), .out(n339) );
  aoi22 U530 ( .a(current_floor_elevator1[55]), .b(n312), .c(
        current_floor_output_elevator1[55]), .d(n313), .out(n338) );
  nand2 U531 ( .a(n340), .b(n341), .out(n911) );
  aoi22 U532 ( .a(n177), .b(N99), .c(N101), .d(n311), .out(n341) );
  aoi22 U533 ( .a(current_floor_elevator1[54]), .b(n312), .c(
        current_floor_output_elevator1[54]), .d(n313), .out(n340) );
  nand2 U534 ( .a(n342), .b(n343), .out(n912) );
  aoi22 U535 ( .a(n177), .b(N100), .c(N102), .d(n311), .out(n343) );
  aoi22 U536 ( .a(current_floor_elevator1[53]), .b(n312), .c(
        current_floor_output_elevator1[53]), .d(n313), .out(n342) );
  nand2 U537 ( .a(n344), .b(n345), .out(n913) );
  aoi22 U538 ( .a(n177), .b(N101), .c(N103), .d(n311), .out(n345) );
  aoi22 U539 ( .a(current_floor_elevator1[52]), .b(n312), .c(
        current_floor_output_elevator1[52]), .d(n313), .out(n344) );
  nand2 U540 ( .a(n346), .b(n347), .out(n914) );
  aoi22 U541 ( .a(n177), .b(N102), .c(N104), .d(n311), .out(n347) );
  aoi22 U542 ( .a(current_floor_elevator1[51]), .b(n312), .c(
        current_floor_output_elevator1[51]), .d(n313), .out(n346) );
  nand2 U543 ( .a(n348), .b(n349), .out(n915) );
  aoi22 U544 ( .a(n177), .b(N103), .c(N105), .d(n311), .out(n349) );
  aoi22 U545 ( .a(current_floor_elevator1[50]), .b(n312), .c(
        current_floor_output_elevator1[50]), .d(n313), .out(n348) );
  nand2 U546 ( .a(n350), .b(n351), .out(n961) );
  aoi22 U547 ( .a(n177), .b(N149), .c(N151), .d(n311), .out(n351) );
  aoi22 U548 ( .a(current_floor_elevator1[4]), .b(n312), .c(
        current_floor_output_elevator1[4]), .d(n313), .out(n350) );
  nand2 U549 ( .a(n352), .b(n353), .out(n916) );
  aoi22 U550 ( .a(n177), .b(N104), .c(N106), .d(n311), .out(n353) );
  aoi22 U551 ( .a(current_floor_elevator1[49]), .b(n312), .c(
        current_floor_output_elevator1[49]), .d(n313), .out(n352) );
  nand2 U552 ( .a(n354), .b(n355), .out(n917) );
  aoi22 U553 ( .a(n177), .b(N105), .c(N107), .d(n311), .out(n355) );
  aoi22 U554 ( .a(current_floor_elevator1[48]), .b(n312), .c(
        current_floor_output_elevator1[48]), .d(n313), .out(n354) );
  nand2 U555 ( .a(n356), .b(n357), .out(n918) );
  aoi22 U556 ( .a(n177), .b(N106), .c(N108), .d(n311), .out(n357) );
  aoi22 U557 ( .a(current_floor_elevator1[47]), .b(n312), .c(
        current_floor_output_elevator1[47]), .d(n313), .out(n356) );
  nand2 U558 ( .a(n358), .b(n359), .out(n919) );
  aoi22 U559 ( .a(n177), .b(N107), .c(N109), .d(n311), .out(n359) );
  aoi22 U560 ( .a(current_floor_elevator1[46]), .b(n312), .c(
        current_floor_output_elevator1[46]), .d(n313), .out(n358) );
  nand2 U561 ( .a(n360), .b(n361), .out(n920) );
  aoi22 U562 ( .a(n177), .b(N108), .c(N110), .d(n311), .out(n361) );
  aoi22 U563 ( .a(current_floor_elevator1[45]), .b(n312), .c(
        current_floor_output_elevator1[45]), .d(n313), .out(n360) );
  nand2 U564 ( .a(n362), .b(n363), .out(n921) );
  aoi22 U565 ( .a(n177), .b(N109), .c(N111), .d(n311), .out(n363) );
  aoi22 U566 ( .a(current_floor_elevator1[44]), .b(n312), .c(
        current_floor_output_elevator1[44]), .d(n313), .out(n362) );
  nand2 U567 ( .a(n364), .b(n365), .out(n922) );
  aoi22 U568 ( .a(n177), .b(N110), .c(N112), .d(n311), .out(n365) );
  aoi22 U569 ( .a(current_floor_elevator1[43]), .b(n312), .c(
        current_floor_output_elevator1[43]), .d(n313), .out(n364) );
  nand2 U570 ( .a(n366), .b(n367), .out(n923) );
  aoi22 U571 ( .a(n177), .b(N111), .c(N113), .d(n311), .out(n367) );
  aoi22 U572 ( .a(current_floor_elevator1[42]), .b(n312), .c(
        current_floor_output_elevator1[42]), .d(n313), .out(n366) );
  nand2 U573 ( .a(n368), .b(n369), .out(n924) );
  aoi22 U574 ( .a(n177), .b(N112), .c(N114), .d(n311), .out(n369) );
  aoi22 U575 ( .a(current_floor_elevator1[41]), .b(n312), .c(
        current_floor_output_elevator1[41]), .d(n313), .out(n368) );
  nand2 U576 ( .a(n370), .b(n371), .out(n925) );
  aoi22 U577 ( .a(n177), .b(N113), .c(N115), .d(n311), .out(n371) );
  aoi22 U578 ( .a(current_floor_elevator1[40]), .b(n312), .c(
        current_floor_output_elevator1[40]), .d(n313), .out(n370) );
  nand2 U579 ( .a(n372), .b(n373), .out(n962) );
  aoi22 U580 ( .a(n177), .b(N150), .c(N152), .d(n311), .out(n373) );
  aoi22 U581 ( .a(current_floor_elevator1[3]), .b(n312), .c(
        current_floor_output_elevator1[3]), .d(n313), .out(n372) );
  nand2 U582 ( .a(n374), .b(n375), .out(n926) );
  aoi22 U583 ( .a(n177), .b(N114), .c(N116), .d(n311), .out(n375) );
  aoi22 U584 ( .a(current_floor_elevator1[39]), .b(n312), .c(
        current_floor_output_elevator1[39]), .d(n313), .out(n374) );
  nand2 U585 ( .a(n376), .b(n377), .out(n927) );
  aoi22 U586 ( .a(n177), .b(N115), .c(N117), .d(n311), .out(n377) );
  aoi22 U587 ( .a(current_floor_elevator1[38]), .b(n312), .c(
        current_floor_output_elevator1[38]), .d(n313), .out(n376) );
  nand2 U588 ( .a(n378), .b(n379), .out(n928) );
  aoi22 U589 ( .a(n177), .b(N116), .c(N118), .d(n311), .out(n379) );
  aoi22 U590 ( .a(current_floor_elevator1[37]), .b(n312), .c(
        current_floor_output_elevator1[37]), .d(n313), .out(n378) );
  nand2 U591 ( .a(n380), .b(n381), .out(n929) );
  aoi22 U592 ( .a(n177), .b(N117), .c(N119), .d(n311), .out(n381) );
  aoi22 U593 ( .a(current_floor_elevator1[36]), .b(n312), .c(
        current_floor_output_elevator1[36]), .d(n313), .out(n380) );
  nand2 U594 ( .a(n382), .b(n383), .out(n930) );
  aoi22 U595 ( .a(n177), .b(N118), .c(N120), .d(n311), .out(n383) );
  aoi22 U596 ( .a(current_floor_elevator1[35]), .b(n312), .c(
        current_floor_output_elevator1[35]), .d(n313), .out(n382) );
  nand2 U597 ( .a(n384), .b(n385), .out(n931) );
  aoi22 U598 ( .a(n177), .b(N119), .c(N121), .d(n311), .out(n385) );
  aoi22 U599 ( .a(current_floor_elevator1[34]), .b(n312), .c(
        current_floor_output_elevator1[34]), .d(n313), .out(n384) );
  nand2 U600 ( .a(n386), .b(n387), .out(n932) );
  aoi22 U601 ( .a(n177), .b(N120), .c(N122), .d(n311), .out(n387) );
  aoi22 U602 ( .a(current_floor_elevator1[33]), .b(n312), .c(
        current_floor_output_elevator1[33]), .d(n313), .out(n386) );
  nand2 U603 ( .a(n388), .b(n389), .out(n933) );
  aoi22 U604 ( .a(n177), .b(N121), .c(N123), .d(n311), .out(n389) );
  aoi22 U605 ( .a(current_floor_elevator1[32]), .b(n312), .c(
        current_floor_output_elevator1[32]), .d(n313), .out(n388) );
  nand2 U606 ( .a(n390), .b(n391), .out(n934) );
  aoi22 U607 ( .a(n177), .b(N122), .c(N124), .d(n311), .out(n391) );
  aoi22 U608 ( .a(current_floor_elevator1[31]), .b(n312), .c(
        current_floor_output_elevator1[31]), .d(n313), .out(n390) );
  nand2 U609 ( .a(n392), .b(n393), .out(n935) );
  aoi22 U610 ( .a(n177), .b(N123), .c(N125), .d(n311), .out(n393) );
  aoi22 U611 ( .a(current_floor_elevator1[30]), .b(n312), .c(
        current_floor_output_elevator1[30]), .d(n313), .out(n392) );
  nand2 U612 ( .a(n394), .b(n395), .out(n963) );
  aoi22 U613 ( .a(n177), .b(N151), .c(N153), .d(n311), .out(n395) );
  aoi22 U614 ( .a(current_floor_elevator1[2]), .b(n312), .c(
        current_floor_output_elevator1[2]), .d(n313), .out(n394) );
  nand2 U615 ( .a(n396), .b(n397), .out(n936) );
  aoi22 U616 ( .a(n177), .b(N124), .c(N126), .d(n311), .out(n397) );
  aoi22 U617 ( .a(current_floor_elevator1[29]), .b(n312), .c(
        current_floor_output_elevator1[29]), .d(n313), .out(n396) );
  nand2 U618 ( .a(n398), .b(n399), .out(n937) );
  aoi22 U619 ( .a(n177), .b(N125), .c(N127), .d(n311), .out(n399) );
  aoi22 U620 ( .a(current_floor_elevator1[28]), .b(n312), .c(
        current_floor_output_elevator1[28]), .d(n313), .out(n398) );
  nand2 U621 ( .a(n400), .b(n401), .out(n938) );
  aoi22 U622 ( .a(n177), .b(N126), .c(N128), .d(n311), .out(n401) );
  aoi22 U623 ( .a(current_floor_elevator1[27]), .b(n312), .c(
        current_floor_output_elevator1[27]), .d(n313), .out(n400) );
  nand2 U624 ( .a(n402), .b(n403), .out(n939) );
  aoi22 U625 ( .a(n177), .b(N127), .c(N129), .d(n311), .out(n403) );
  aoi22 U626 ( .a(current_floor_elevator1[26]), .b(n312), .c(
        current_floor_output_elevator1[26]), .d(n313), .out(n402) );
  nand2 U627 ( .a(n404), .b(n405), .out(n940) );
  aoi22 U628 ( .a(n177), .b(N128), .c(N130), .d(n311), .out(n405) );
  aoi22 U629 ( .a(current_floor_elevator1[25]), .b(n312), .c(
        current_floor_output_elevator1[25]), .d(n313), .out(n404) );
  nand2 U630 ( .a(n406), .b(n407), .out(n941) );
  aoi22 U631 ( .a(n177), .b(N129), .c(N131), .d(n311), .out(n407) );
  aoi22 U632 ( .a(current_floor_elevator1[24]), .b(n312), .c(
        current_floor_output_elevator1[24]), .d(n313), .out(n406) );
  nand2 U633 ( .a(n408), .b(n409), .out(n942) );
  aoi22 U634 ( .a(n177), .b(N130), .c(N132), .d(n311), .out(n409) );
  aoi22 U635 ( .a(current_floor_elevator1[23]), .b(n312), .c(
        current_floor_output_elevator1[23]), .d(n313), .out(n408) );
  nand2 U636 ( .a(n410), .b(n411), .out(n943) );
  aoi22 U637 ( .a(n177), .b(N131), .c(N133), .d(n311), .out(n411) );
  aoi22 U638 ( .a(current_floor_elevator1[22]), .b(n312), .c(
        current_floor_output_elevator1[22]), .d(n313), .out(n410) );
  nand2 U639 ( .a(n412), .b(n413), .out(n944) );
  aoi22 U640 ( .a(n177), .b(N132), .c(N134), .d(n311), .out(n413) );
  aoi22 U641 ( .a(current_floor_elevator1[21]), .b(n312), .c(
        current_floor_output_elevator1[21]), .d(n313), .out(n412) );
  nand2 U642 ( .a(n414), .b(n415), .out(n945) );
  aoi22 U643 ( .a(n177), .b(N133), .c(N135), .d(n311), .out(n415) );
  aoi22 U644 ( .a(current_floor_elevator1[20]), .b(n312), .c(
        current_floor_output_elevator1[20]), .d(n313), .out(n414) );
  nand2 U645 ( .a(n416), .b(n417), .out(n964) );
  aoi22 U646 ( .a(n177), .b(N152), .c(N154), .d(n311), .out(n417) );
  aoi22 U647 ( .a(current_floor_elevator1[1]), .b(n312), .c(
        current_floor_output_elevator1[1]), .d(n313), .out(n416) );
  nand2 U648 ( .a(n418), .b(n419), .out(n946) );
  aoi22 U649 ( .a(n177), .b(N134), .c(N136), .d(n311), .out(n419) );
  aoi22 U650 ( .a(current_floor_elevator1[19]), .b(n312), .c(
        current_floor_output_elevator1[19]), .d(n313), .out(n418) );
  nand2 U651 ( .a(n420), .b(n421), .out(n947) );
  aoi22 U652 ( .a(n177), .b(N135), .c(N137), .d(n311), .out(n421) );
  aoi22 U653 ( .a(current_floor_elevator1[18]), .b(n312), .c(
        current_floor_output_elevator1[18]), .d(n313), .out(n420) );
  nand2 U654 ( .a(n422), .b(n423), .out(n948) );
  aoi22 U655 ( .a(n177), .b(N136), .c(N138), .d(n311), .out(n423) );
  aoi22 U656 ( .a(current_floor_elevator1[17]), .b(n312), .c(
        current_floor_output_elevator1[17]), .d(n313), .out(n422) );
  nand2 U657 ( .a(n424), .b(n425), .out(n949) );
  aoi22 U658 ( .a(n177), .b(N137), .c(N139), .d(n311), .out(n425) );
  aoi22 U659 ( .a(current_floor_elevator1[16]), .b(n312), .c(
        current_floor_output_elevator1[16]), .d(n313), .out(n424) );
  nand2 U660 ( .a(n426), .b(n427), .out(n950) );
  aoi22 U661 ( .a(n177), .b(N138), .c(N140), .d(n311), .out(n427) );
  aoi22 U662 ( .a(current_floor_elevator1[15]), .b(n312), .c(
        current_floor_output_elevator1[15]), .d(n313), .out(n426) );
  nand2 U663 ( .a(n428), .b(n429), .out(n951) );
  aoi22 U664 ( .a(n177), .b(N139), .c(N141), .d(n311), .out(n429) );
  aoi22 U665 ( .a(current_floor_elevator1[14]), .b(n312), .c(
        current_floor_output_elevator1[14]), .d(n313), .out(n428) );
  nand2 U666 ( .a(n430), .b(n431), .out(n952) );
  aoi22 U667 ( .a(n177), .b(N140), .c(N142), .d(n311), .out(n431) );
  aoi22 U668 ( .a(current_floor_elevator1[13]), .b(n312), .c(
        current_floor_output_elevator1[13]), .d(n313), .out(n430) );
  nand2 U669 ( .a(n432), .b(n433), .out(n953) );
  aoi22 U670 ( .a(n177), .b(N141), .c(N143), .d(n311), .out(n433) );
  aoi22 U671 ( .a(current_floor_elevator1[12]), .b(n312), .c(
        current_floor_output_elevator1[12]), .d(n313), .out(n432) );
  nand2 U672 ( .a(n434), .b(n435), .out(n954) );
  aoi22 U673 ( .a(n177), .b(N142), .c(N144), .d(n311), .out(n435) );
  aoi22 U674 ( .a(current_floor_elevator1[11]), .b(n312), .c(
        current_floor_output_elevator1[11]), .d(n313), .out(n434) );
  nand2 U675 ( .a(n436), .b(n437), .out(n955) );
  aoi22 U676 ( .a(n177), .b(N143), .c(N145), .d(n311), .out(n437) );
  aoi22 U677 ( .a(current_floor_elevator1[10]), .b(n312), .c(
        current_floor_output_elevator1[10]), .d(n313), .out(n436) );
  nand2 U678 ( .a(n438), .b(n439), .out(n965) );
  nand2 U679 ( .a(current_floor_output_elevator1[0]), .b(n313), .out(n439) );
  aoi22 U680 ( .a(n177), .b(N153), .c(current_floor_elevator1[0]), .d(n312), 
        .out(n438) );
  nor2 U681 ( .a(n313), .b(n1172), .out(n312) );
  nand3 U682 ( .a(n440), .b(n32), .c(n441), .out(n967) );
  nand2 U683 ( .a(in_emergency_elevator2), .b(n28), .out(n441) );
  nand2 U684 ( .a(N509), .b(n28), .out(n32) );
  inv U685 ( .in(n1170), .out(n28) );
  nand3 U686 ( .a(n182), .b(n1169), .c(arrived_elevator2), .out(n440) );
  nor3 U687 ( .a(n180), .b(n1595), .c(n172), .out(n182) );
  nor2 U688 ( .a(n180), .b(n1167), .out(n172) );
  nand2 U689 ( .a(N507), .b(n1169), .out(n1167) );
  inv U690 ( .in(n1168), .out(n180) );
  nand2 U691 ( .a(N505), .b(n1169), .out(n1168) );
  inv U692 ( .in(in_emergency_elevator2), .out(n1169) );
  nand3 U694 ( .a(n442), .b(n167), .c(n443), .out(n899) );
  nand2 U695 ( .a(in_emergency_elevator1), .b(n444), .out(n443) );
  nand2 U696 ( .a(N225), .b(n444), .out(n167) );
  inv U697 ( .in(n1172), .out(n444) );
  nand3 U698 ( .a(n313), .b(n1171), .c(arrived_elevator1), .out(n442) );
  nor3 U699 ( .a(n311), .b(n1640), .c(n177), .out(n313) );
  nor2 U700 ( .a(n311), .b(n1165), .out(n177) );
  nand2 U701 ( .a(N223), .b(n1171), .out(n1165) );
  inv U702 ( .in(n1166), .out(n311) );
  nand2 U703 ( .a(N221), .b(n1171), .out(n1166) );
  inv U704 ( .in(in_emergency_elevator1), .out(n1171) );
  nand2 U705 ( .a(n881), .b(n880), .out(N99) );
  nand2 U706 ( .a(n883), .b(n882), .out(N98) );
  nand2 U707 ( .a(n885), .b(n884), .out(N97) );
  nand2 U708 ( .a(n887), .b(n886), .out(N96) );
  nand2 U709 ( .a(n889), .b(n888), .out(N95) );
  nand2 U710 ( .a(n891), .b(n890), .out(N94) );
  nand2 U711 ( .a(n893), .b(n892), .out(N93) );
  nand2 U712 ( .a(n895), .b(n894), .out(N92) );
  nand2 U713 ( .a(n897), .b(n896), .out(\r125/SB ) );
  oai12 U714 ( .b(n1640), .c(n445), .a(n446), .out(N90) );
  nand2 U715 ( .a(\eq_42_3/SB ), .b(n1640), .out(n446) );
  oai12 U716 ( .b(n1640), .c(n447), .a(n448), .out(N89) );
  nand2 U717 ( .a(destination_floor_elevator1[62]), .b(n1640), .out(n448) );
  oai12 U718 ( .b(n1640), .c(n449), .a(n450), .out(N88) );
  nand2 U719 ( .a(destination_floor_elevator1[61]), .b(n1640), .out(n450) );
  oai12 U720 ( .b(n1640), .c(n451), .a(n452), .out(N87) );
  nand2 U721 ( .a(destination_floor_elevator1[60]), .b(n1640), .out(n452) );
  oai12 U722 ( .b(n1640), .c(n453), .a(n454), .out(N86) );
  nand2 U723 ( .a(destination_floor_elevator1[59]), .b(n1641), .out(n454) );
  oai12 U724 ( .b(n1641), .c(n455), .a(n456), .out(N85) );
  nand2 U725 ( .a(destination_floor_elevator1[58]), .b(n1641), .out(n456) );
  oai12 U726 ( .b(n1641), .c(n457), .a(n458), .out(N84) );
  nand2 U727 ( .a(destination_floor_elevator1[57]), .b(n1641), .out(n458) );
  oai12 U728 ( .b(n1641), .c(n459), .a(n460), .out(N83) );
  nand2 U729 ( .a(destination_floor_elevator1[56]), .b(n1641), .out(n460) );
  oai12 U730 ( .b(n1641), .c(n461), .a(n462), .out(N82) );
  nand2 U731 ( .a(destination_floor_elevator1[55]), .b(n1641), .out(n462) );
  oai12 U732 ( .b(n1641), .c(n463), .a(n464), .out(N81) );
  nand2 U733 ( .a(destination_floor_elevator1[54]), .b(n1641), .out(n464) );
  oai12 U734 ( .b(n1641), .c(n465), .a(n466), .out(N80) );
  nand2 U735 ( .a(destination_floor_elevator1[53]), .b(n1642), .out(n466) );
  oai12 U736 ( .b(n1642), .c(n467), .a(n468), .out(N79) );
  nand2 U737 ( .a(destination_floor_elevator1[52]), .b(n1642), .out(n468) );
  oai12 U738 ( .b(n1642), .c(n469), .a(n470), .out(N78) );
  nand2 U739 ( .a(destination_floor_elevator1[51]), .b(n1642), .out(n470) );
  oai12 U740 ( .b(n1642), .c(n471), .a(n472), .out(N77) );
  nand2 U741 ( .a(destination_floor_elevator1[50]), .b(n1642), .out(n472) );
  nand2 U742 ( .a(n1662), .b(n473), .out(N76) );
  oai12 U744 ( .b(n1642), .c(n474), .a(n475), .out(N75) );
  nand2 U745 ( .a(destination_floor_elevator1[49]), .b(n1642), .out(n475) );
  oai12 U746 ( .b(n1642), .c(n476), .a(n477), .out(N74) );
  nand2 U747 ( .a(destination_floor_elevator1[48]), .b(n1642), .out(n477) );
  oai12 U748 ( .b(n1642), .c(n478), .a(n479), .out(N73) );
  nand2 U749 ( .a(destination_floor_elevator1[47]), .b(n1643), .out(n479) );
  oai12 U750 ( .b(n1643), .c(n480), .a(n481), .out(N72) );
  nand2 U751 ( .a(destination_floor_elevator1[46]), .b(n1643), .out(n481) );
  oai12 U752 ( .b(n1643), .c(n482), .a(n483), .out(N71) );
  nand2 U753 ( .a(destination_floor_elevator1[45]), .b(n1643), .out(n483) );
  oai12 U754 ( .b(n1643), .c(n484), .a(n485), .out(N70) );
  nand2 U755 ( .a(destination_floor_elevator1[44]), .b(n1643), .out(n485) );
  oai12 U756 ( .b(n1643), .c(n486), .a(n487), .out(N69) );
  nand2 U757 ( .a(destination_floor_elevator1[43]), .b(n1643), .out(n487) );
  oai12 U758 ( .b(n1643), .c(n488), .a(n489), .out(N68) );
  nand2 U759 ( .a(destination_floor_elevator1[42]), .b(n1643), .out(n489) );
  oai12 U760 ( .b(n1643), .c(n490), .a(n491), .out(N67) );
  nand2 U761 ( .a(destination_floor_elevator1[41]), .b(n1644), .out(n491) );
  oai12 U762 ( .b(n1644), .c(n492), .a(n493), .out(N66) );
  nand2 U763 ( .a(destination_floor_elevator1[40]), .b(n1644), .out(n493) );
  oai12 U764 ( .b(n1644), .c(n494), .a(n495), .out(N65) );
  nand2 U765 ( .a(destination_floor_elevator1[39]), .b(n1644), .out(n495) );
  oai12 U766 ( .b(n1644), .c(n496), .a(n497), .out(N64) );
  nand2 U767 ( .a(destination_floor_elevator1[38]), .b(n1644), .out(n497) );
  oai12 U768 ( .b(n1644), .c(n498), .a(n499), .out(N63) );
  nand2 U769 ( .a(destination_floor_elevator1[37]), .b(n1644), .out(n499) );
  oai12 U770 ( .b(n1644), .c(n500), .a(n501), .out(N62) );
  nand2 U771 ( .a(destination_floor_elevator1[36]), .b(n1644), .out(n501) );
  oai12 U772 ( .b(n1644), .c(n502), .a(n503), .out(N61) );
  nand2 U773 ( .a(destination_floor_elevator1[35]), .b(n1645), .out(n503) );
  oai12 U774 ( .b(n1645), .c(n504), .a(n505), .out(N60) );
  nand2 U775 ( .a(destination_floor_elevator1[34]), .b(n1645), .out(n505) );
  oai12 U776 ( .b(n1645), .c(n506), .a(n507), .out(N59) );
  nand2 U777 ( .a(destination_floor_elevator1[33]), .b(n1645), .out(n507) );
  oai12 U778 ( .b(n1645), .c(n508), .a(n509), .out(N58) );
  nand2 U779 ( .a(destination_floor_elevator1[32]), .b(n1645), .out(n509) );
  oai12 U780 ( .b(n1645), .c(n510), .a(n511), .out(N57) );
  nand2 U781 ( .a(destination_floor_elevator1[31]), .b(n1645), .out(n511) );
  oai12 U782 ( .b(n1645), .c(n512), .a(n513), .out(N56) );
  nand2 U783 ( .a(destination_floor_elevator1[30]), .b(n1645), .out(n513) );
  oai12 U784 ( .b(n1645), .c(n514), .a(n515), .out(N55) );
  nand2 U785 ( .a(destination_floor_elevator1[29]), .b(n1646), .out(n515) );
  oai12 U786 ( .b(n1646), .c(n516), .a(n517), .out(N54) );
  nand2 U787 ( .a(destination_floor_elevator1[28]), .b(n1646), .out(n517) );
  oai12 U788 ( .b(n1646), .c(n518), .a(n519), .out(N53) );
  nand2 U789 ( .a(destination_floor_elevator1[27]), .b(n1646), .out(n519) );
  oai12 U790 ( .b(n1646), .c(n520), .a(n521), .out(N52) );
  nand2 U791 ( .a(destination_floor_elevator1[26]), .b(n1646), .out(n521) );
  oai12 U792 ( .b(n1646), .c(n522), .a(n523), .out(N51) );
  nand2 U793 ( .a(destination_floor_elevator1[25]), .b(n1646), .out(n523) );
  oai12 U794 ( .b(n1646), .c(n524), .a(n525), .out(N50) );
  nand2 U795 ( .a(destination_floor_elevator1[24]), .b(n1646), .out(n525) );
  oai12 U796 ( .b(n1646), .c(n526), .a(n527), .out(N49) );
  nand2 U797 ( .a(destination_floor_elevator1[23]), .b(n1647), .out(n527) );
  oai12 U798 ( .b(n1647), .c(n528), .a(n529), .out(N48) );
  nand2 U799 ( .a(destination_floor_elevator1[22]), .b(n1647), .out(n529) );
  oai12 U800 ( .b(n1647), .c(n530), .a(n531), .out(N47) );
  nand2 U801 ( .a(destination_floor_elevator1[21]), .b(n1647), .out(n531) );
  oai12 U802 ( .b(n1647), .c(n532), .a(n533), .out(N46) );
  nand2 U803 ( .a(destination_floor_elevator1[20]), .b(n1647), .out(n533) );
  oai12 U804 ( .b(n1647), .c(n534), .a(n535), .out(N45) );
  nand2 U805 ( .a(destination_floor_elevator1[19]), .b(n1647), .out(n535) );
  oai12 U806 ( .b(n1647), .c(n536), .a(n537), .out(N44) );
  nand2 U807 ( .a(destination_floor_elevator1[18]), .b(n1647), .out(n537) );
  nand2 U808 ( .a(n647), .b(n646), .out(N438) );
  nand2 U809 ( .a(n643), .b(n642), .out(N437) );
  nand2 U810 ( .a(n645), .b(n644), .out(N436) );
  nand2 U811 ( .a(n649), .b(n648), .out(N435) );
  nand2 U812 ( .a(n651), .b(n650), .out(N434) );
  nand2 U813 ( .a(n653), .b(n652), .out(N433) );
  nand2 U814 ( .a(n655), .b(n654), .out(N432) );
  nand2 U815 ( .a(n657), .b(n656), .out(N431) );
  nand2 U816 ( .a(n659), .b(n658), .out(N430) );
  oai12 U817 ( .b(n1647), .c(n538), .a(n539), .out(N43) );
  nand2 U818 ( .a(destination_floor_elevator1[17]), .b(n1648), .out(n539) );
  nand2 U819 ( .a(n661), .b(n660), .out(N429) );
  nand2 U820 ( .a(n663), .b(n662), .out(N428) );
  nand2 U821 ( .a(n665), .b(n664), .out(N427) );
  nand2 U822 ( .a(n667), .b(n666), .out(N426) );
  nand2 U823 ( .a(n669), .b(n668), .out(N425) );
  nand2 U824 ( .a(n671), .b(n670), .out(N424) );
  nand2 U825 ( .a(n673), .b(n672), .out(N423) );
  nand2 U826 ( .a(n675), .b(n674), .out(N422) );
  nand2 U827 ( .a(n677), .b(n676), .out(N421) );
  nand2 U828 ( .a(n679), .b(n678), .out(N420) );
  oai12 U829 ( .b(n1648), .c(n540), .a(n541), .out(N42) );
  nand2 U830 ( .a(destination_floor_elevator1[16]), .b(n1648), .out(n541) );
  nand2 U831 ( .a(n681), .b(n680), .out(N419) );
  nand2 U832 ( .a(n683), .b(n682), .out(N418) );
  nand2 U833 ( .a(n685), .b(n684), .out(N417) );
  nand2 U834 ( .a(n687), .b(n686), .out(N416) );
  nand2 U835 ( .a(n689), .b(n688), .out(N415) );
  nand2 U836 ( .a(n691), .b(n690), .out(N414) );
  nand2 U837 ( .a(n693), .b(n692), .out(N413) );
  nand2 U838 ( .a(n695), .b(n694), .out(N412) );
  nand2 U839 ( .a(n697), .b(n696), .out(N411) );
  nand2 U840 ( .a(n699), .b(n698), .out(N410) );
  oai12 U841 ( .b(n1648), .c(n542), .a(n543), .out(N41) );
  nand2 U842 ( .a(destination_floor_elevator1[15]), .b(n1648), .out(n543) );
  nand2 U843 ( .a(n701), .b(n700), .out(N409) );
  nand2 U844 ( .a(n703), .b(n702), .out(N408) );
  nand2 U845 ( .a(n705), .b(n704), .out(N407) );
  nand2 U846 ( .a(n707), .b(n706), .out(N406) );
  nand2 U847 ( .a(n709), .b(n708), .out(N405) );
  nand2 U848 ( .a(n711), .b(n710), .out(N404) );
  nand2 U849 ( .a(n713), .b(n712), .out(N403) );
  nand2 U850 ( .a(n715), .b(n714), .out(N402) );
  nand2 U851 ( .a(n717), .b(n716), .out(N401) );
  nand2 U852 ( .a(n719), .b(n718), .out(N400) );
  oai12 U853 ( .b(n1648), .c(n544), .a(n545), .out(N40) );
  nand2 U854 ( .a(destination_floor_elevator1[14]), .b(n1648), .out(n545) );
  nand2 U855 ( .a(n721), .b(n720), .out(N399) );
  nand2 U856 ( .a(n723), .b(n722), .out(N398) );
  nand2 U857 ( .a(n725), .b(n724), .out(N397) );
  nand2 U858 ( .a(n727), .b(n726), .out(N396) );
  nand2 U859 ( .a(n729), .b(n728), .out(N395) );
  nand2 U860 ( .a(n731), .b(n730), .out(N394) );
  nand2 U861 ( .a(n733), .b(n732), .out(N393) );
  nand2 U862 ( .a(n735), .b(n734), .out(N392) );
  nand2 U863 ( .a(n737), .b(n736), .out(N391) );
  nand2 U864 ( .a(n739), .b(n738), .out(N390) );
  oai12 U865 ( .b(n1648), .c(n546), .a(n547), .out(N39) );
  nand2 U866 ( .a(destination_floor_elevator1[13]), .b(n1648), .out(n547) );
  nand2 U867 ( .a(n741), .b(n740), .out(N389) );
  nand2 U868 ( .a(n743), .b(n742), .out(N388) );
  nand2 U869 ( .a(n745), .b(n744), .out(N387) );
  nand2 U870 ( .a(n747), .b(n746), .out(N386) );
  nand2 U871 ( .a(n749), .b(n748), .out(N385) );
  nand2 U872 ( .a(n751), .b(n750), .out(N384) );
  nand2 U873 ( .a(n753), .b(n752), .out(N383) );
  nand2 U874 ( .a(n755), .b(n754), .out(N382) );
  nand2 U875 ( .a(n757), .b(n756), .out(N381) );
  nand2 U876 ( .a(n759), .b(n758), .out(N380) );
  oai12 U877 ( .b(n1648), .c(n548), .a(n549), .out(N38) );
  nand2 U878 ( .a(destination_floor_elevator1[12]), .b(n1648), .out(n549) );
  nand2 U879 ( .a(n761), .b(n760), .out(N379) );
  nand2 U880 ( .a(n763), .b(n762), .out(N378) );
  nand2 U881 ( .a(n765), .b(n764), .out(N377) );
  nand2 U882 ( .a(n767), .b(n766), .out(N376) );
  nand2 U883 ( .a(n769), .b(n768), .out(\r126/SB ) );
  oai12 U884 ( .b(n1595), .c(n445), .a(n550), .out(N374) );
  nand2 U885 ( .a(\eq_47_3/SB ), .b(n1595), .out(n550) );
  inv U886 ( .in(\ne_47/SB ), .out(n445) );
  oai12 U887 ( .b(n1595), .c(n447), .a(n551), .out(N373) );
  nand2 U888 ( .a(destination_floor_elevator2[62]), .b(n1595), .out(n551) );
  inv U889 ( .in(requested_floor[62]), .out(n447) );
  oai12 U890 ( .b(n1595), .c(n449), .a(n552), .out(N372) );
  nand2 U891 ( .a(destination_floor_elevator2[61]), .b(n1595), .out(n552) );
  inv U892 ( .in(requested_floor[61]), .out(n449) );
  oai12 U893 ( .b(n1595), .c(n451), .a(n553), .out(N371) );
  nand2 U894 ( .a(destination_floor_elevator2[60]), .b(n1595), .out(n553) );
  inv U895 ( .in(requested_floor[60]), .out(n451) );
  oai12 U896 ( .b(n1595), .c(n453), .a(n554), .out(N370) );
  nand2 U897 ( .a(destination_floor_elevator2[59]), .b(n1596), .out(n554) );
  inv U898 ( .in(requested_floor[59]), .out(n453) );
  oai12 U899 ( .b(n1648), .c(n555), .a(n556), .out(N37) );
  nand2 U900 ( .a(destination_floor_elevator1[11]), .b(n1649), .out(n556) );
  oai12 U901 ( .b(n1596), .c(n455), .a(n557), .out(N369) );
  nand2 U902 ( .a(destination_floor_elevator2[58]), .b(n1596), .out(n557) );
  inv U903 ( .in(requested_floor[58]), .out(n455) );
  oai12 U904 ( .b(n1596), .c(n457), .a(n558), .out(N368) );
  nand2 U905 ( .a(destination_floor_elevator2[57]), .b(n1596), .out(n558) );
  inv U906 ( .in(requested_floor[57]), .out(n457) );
  oai12 U907 ( .b(n1596), .c(n459), .a(n559), .out(N367) );
  nand2 U908 ( .a(destination_floor_elevator2[56]), .b(n1596), .out(n559) );
  inv U909 ( .in(requested_floor[56]), .out(n459) );
  oai12 U910 ( .b(n1596), .c(n461), .a(n560), .out(N366) );
  nand2 U911 ( .a(destination_floor_elevator2[55]), .b(n1596), .out(n560) );
  inv U912 ( .in(requested_floor[55]), .out(n461) );
  oai12 U913 ( .b(n1596), .c(n463), .a(n561), .out(N365) );
  nand2 U914 ( .a(destination_floor_elevator2[54]), .b(n1596), .out(n561) );
  inv U915 ( .in(requested_floor[54]), .out(n463) );
  oai12 U916 ( .b(n1596), .c(n465), .a(n562), .out(N364) );
  nand2 U917 ( .a(destination_floor_elevator2[53]), .b(n1597), .out(n562) );
  inv U918 ( .in(requested_floor[53]), .out(n465) );
  oai12 U919 ( .b(n1597), .c(n467), .a(n563), .out(N363) );
  nand2 U920 ( .a(destination_floor_elevator2[52]), .b(n1597), .out(n563) );
  inv U921 ( .in(requested_floor[52]), .out(n467) );
  oai12 U922 ( .b(n1597), .c(n469), .a(n564), .out(N362) );
  nand2 U923 ( .a(destination_floor_elevator2[51]), .b(n1597), .out(n564) );
  inv U924 ( .in(requested_floor[51]), .out(n469) );
  oai12 U925 ( .b(n1597), .c(n471), .a(n565), .out(N361) );
  nand2 U926 ( .a(destination_floor_elevator2[50]), .b(n1597), .out(n565) );
  inv U927 ( .in(requested_floor[50]), .out(n471) );
  nand2 U928 ( .a(n1617), .b(n566), .out(N360) );
  nand3 U929 ( .a(n473), .b(n34), .c(N16), .out(n566) );
  inv U930 ( .in(n640), .out(n34) );
  nand2 U931 ( .a(N13), .b(n567), .out(n473) );
  inv U932 ( .in(n641), .out(n567) );
  oai12 U934 ( .b(n1649), .c(n568), .a(n569), .out(N36) );
  nand2 U935 ( .a(destination_floor_elevator1[10]), .b(n1649), .out(n569) );
  oai12 U936 ( .b(n1597), .c(n474), .a(n570), .out(N359) );
  nand2 U937 ( .a(destination_floor_elevator2[49]), .b(n1597), .out(n570) );
  inv U938 ( .in(requested_floor[49]), .out(n474) );
  oai12 U939 ( .b(n1597), .c(n476), .a(n571), .out(N358) );
  nand2 U940 ( .a(destination_floor_elevator2[48]), .b(n1597), .out(n571) );
  inv U941 ( .in(requested_floor[48]), .out(n476) );
  oai12 U942 ( .b(n1597), .c(n478), .a(n572), .out(N357) );
  nand2 U943 ( .a(destination_floor_elevator2[47]), .b(n1598), .out(n572) );
  inv U944 ( .in(requested_floor[47]), .out(n478) );
  oai12 U945 ( .b(n1598), .c(n480), .a(n573), .out(N356) );
  nand2 U946 ( .a(destination_floor_elevator2[46]), .b(n1598), .out(n573) );
  inv U947 ( .in(requested_floor[46]), .out(n480) );
  oai12 U948 ( .b(n1598), .c(n482), .a(n574), .out(N355) );
  nand2 U949 ( .a(destination_floor_elevator2[45]), .b(n1598), .out(n574) );
  inv U950 ( .in(requested_floor[45]), .out(n482) );
  oai12 U951 ( .b(n1598), .c(n484), .a(n575), .out(N354) );
  nand2 U952 ( .a(destination_floor_elevator2[44]), .b(n1598), .out(n575) );
  inv U953 ( .in(requested_floor[44]), .out(n484) );
  oai12 U954 ( .b(n1598), .c(n486), .a(n576), .out(N353) );
  nand2 U955 ( .a(destination_floor_elevator2[43]), .b(n1598), .out(n576) );
  inv U956 ( .in(requested_floor[43]), .out(n486) );
  oai12 U957 ( .b(n1598), .c(n488), .a(n577), .out(N352) );
  nand2 U958 ( .a(destination_floor_elevator2[42]), .b(n1598), .out(n577) );
  inv U959 ( .in(requested_floor[42]), .out(n488) );
  oai12 U960 ( .b(n1598), .c(n490), .a(n578), .out(N351) );
  nand2 U961 ( .a(destination_floor_elevator2[41]), .b(n1599), .out(n578) );
  inv U962 ( .in(requested_floor[41]), .out(n490) );
  oai12 U963 ( .b(n1599), .c(n492), .a(n579), .out(N350) );
  nand2 U964 ( .a(destination_floor_elevator2[40]), .b(n1599), .out(n579) );
  inv U965 ( .in(requested_floor[40]), .out(n492) );
  oai12 U966 ( .b(n1649), .c(n580), .a(n581), .out(N35) );
  nand2 U967 ( .a(n1649), .b(destination_floor_elevator1[9]), .out(n581) );
  oai12 U968 ( .b(n1599), .c(n494), .a(n582), .out(N349) );
  nand2 U969 ( .a(destination_floor_elevator2[39]), .b(n1599), .out(n582) );
  inv U970 ( .in(requested_floor[39]), .out(n494) );
  oai12 U971 ( .b(n1599), .c(n496), .a(n583), .out(N348) );
  nand2 U972 ( .a(destination_floor_elevator2[38]), .b(n1599), .out(n583) );
  inv U973 ( .in(requested_floor[38]), .out(n496) );
  oai12 U974 ( .b(n1599), .c(n498), .a(n584), .out(N347) );
  nand2 U975 ( .a(destination_floor_elevator2[37]), .b(n1599), .out(n584) );
  inv U976 ( .in(requested_floor[37]), .out(n498) );
  oai12 U977 ( .b(n1599), .c(n500), .a(n585), .out(N346) );
  nand2 U978 ( .a(destination_floor_elevator2[36]), .b(n1599), .out(n585) );
  inv U979 ( .in(requested_floor[36]), .out(n500) );
  oai12 U980 ( .b(n1599), .c(n502), .a(n586), .out(N345) );
  nand2 U981 ( .a(destination_floor_elevator2[35]), .b(n1600), .out(n586) );
  inv U982 ( .in(requested_floor[35]), .out(n502) );
  oai12 U983 ( .b(n1600), .c(n504), .a(n587), .out(N344) );
  nand2 U984 ( .a(destination_floor_elevator2[34]), .b(n1600), .out(n587) );
  inv U985 ( .in(requested_floor[34]), .out(n504) );
  oai12 U986 ( .b(n1600), .c(n506), .a(n588), .out(N343) );
  nand2 U987 ( .a(destination_floor_elevator2[33]), .b(n1600), .out(n588) );
  inv U988 ( .in(requested_floor[33]), .out(n506) );
  oai12 U989 ( .b(n1600), .c(n508), .a(n589), .out(N342) );
  nand2 U990 ( .a(destination_floor_elevator2[32]), .b(n1600), .out(n589) );
  inv U991 ( .in(requested_floor[32]), .out(n508) );
  oai12 U992 ( .b(n1600), .c(n510), .a(n590), .out(N341) );
  nand2 U993 ( .a(destination_floor_elevator2[31]), .b(n1600), .out(n590) );
  inv U994 ( .in(requested_floor[31]), .out(n510) );
  oai12 U995 ( .b(n1600), .c(n512), .a(n591), .out(N340) );
  nand2 U996 ( .a(destination_floor_elevator2[30]), .b(n1600), .out(n591) );
  inv U997 ( .in(requested_floor[30]), .out(n512) );
  oai12 U998 ( .b(n1649), .c(n592), .a(n593), .out(N34) );
  nand2 U999 ( .a(destination_floor_elevator1[8]), .b(n1649), .out(n593) );
  oai12 U1000 ( .b(n1600), .c(n514), .a(n594), .out(N339) );
  nand2 U1001 ( .a(destination_floor_elevator2[29]), .b(n1601), .out(n594) );
  inv U1002 ( .in(requested_floor[29]), .out(n514) );
  oai12 U1003 ( .b(n1601), .c(n516), .a(n595), .out(N338) );
  nand2 U1004 ( .a(destination_floor_elevator2[28]), .b(n1601), .out(n595) );
  inv U1005 ( .in(requested_floor[28]), .out(n516) );
  oai12 U1006 ( .b(n1601), .c(n518), .a(n596), .out(N337) );
  nand2 U1007 ( .a(destination_floor_elevator2[27]), .b(n1601), .out(n596) );
  inv U1008 ( .in(requested_floor[27]), .out(n518) );
  oai12 U1009 ( .b(n1601), .c(n520), .a(n597), .out(N336) );
  nand2 U1010 ( .a(destination_floor_elevator2[26]), .b(n1601), .out(n597) );
  inv U1011 ( .in(requested_floor[26]), .out(n520) );
  oai12 U1012 ( .b(n1601), .c(n522), .a(n598), .out(N335) );
  nand2 U1013 ( .a(destination_floor_elevator2[25]), .b(n1601), .out(n598) );
  inv U1014 ( .in(requested_floor[25]), .out(n522) );
  oai12 U1015 ( .b(n1601), .c(n524), .a(n599), .out(N334) );
  nand2 U1016 ( .a(destination_floor_elevator2[24]), .b(n1601), .out(n599) );
  inv U1017 ( .in(requested_floor[24]), .out(n524) );
  oai12 U1018 ( .b(n1601), .c(n526), .a(n600), .out(N333) );
  nand2 U1019 ( .a(destination_floor_elevator2[23]), .b(n1602), .out(n600) );
  inv U1020 ( .in(requested_floor[23]), .out(n526) );
  oai12 U1021 ( .b(n1602), .c(n528), .a(n601), .out(N332) );
  nand2 U1022 ( .a(destination_floor_elevator2[22]), .b(n1602), .out(n601) );
  inv U1023 ( .in(requested_floor[22]), .out(n528) );
  oai12 U1024 ( .b(n1602), .c(n530), .a(n602), .out(N331) );
  nand2 U1025 ( .a(destination_floor_elevator2[21]), .b(n1602), .out(n602) );
  inv U1026 ( .in(requested_floor[21]), .out(n530) );
  oai12 U1027 ( .b(n1602), .c(n532), .a(n603), .out(N330) );
  nand2 U1028 ( .a(destination_floor_elevator2[20]), .b(n1602), .out(n603) );
  inv U1029 ( .in(requested_floor[20]), .out(n532) );
  oai12 U1030 ( .b(n1649), .c(n604), .a(n605), .out(N33) );
  nand2 U1031 ( .a(destination_floor_elevator1[7]), .b(n1649), .out(n605) );
  oai12 U1032 ( .b(n1602), .c(n534), .a(n606), .out(N329) );
  nand2 U1033 ( .a(destination_floor_elevator2[19]), .b(n1602), .out(n606) );
  inv U1034 ( .in(requested_floor[19]), .out(n534) );
  oai12 U1035 ( .b(n1602), .c(n536), .a(n607), .out(N328) );
  nand2 U1036 ( .a(destination_floor_elevator2[18]), .b(n1602), .out(n607) );
  inv U1037 ( .in(requested_floor[18]), .out(n536) );
  oai12 U1038 ( .b(n1602), .c(n538), .a(n608), .out(N327) );
  nand2 U1039 ( .a(destination_floor_elevator2[17]), .b(n1603), .out(n608) );
  inv U1040 ( .in(requested_floor[17]), .out(n538) );
  oai12 U1041 ( .b(n1603), .c(n540), .a(n609), .out(N326) );
  nand2 U1042 ( .a(destination_floor_elevator2[16]), .b(n1603), .out(n609) );
  inv U1043 ( .in(requested_floor[16]), .out(n540) );
  oai12 U1044 ( .b(n1603), .c(n542), .a(n610), .out(N325) );
  nand2 U1045 ( .a(destination_floor_elevator2[15]), .b(n1603), .out(n610) );
  inv U1046 ( .in(requested_floor[15]), .out(n542) );
  oai12 U1047 ( .b(n1603), .c(n544), .a(n611), .out(N324) );
  nand2 U1048 ( .a(destination_floor_elevator2[14]), .b(n1603), .out(n611) );
  inv U1049 ( .in(requested_floor[14]), .out(n544) );
  oai12 U1050 ( .b(n1603), .c(n546), .a(n612), .out(N323) );
  nand2 U1051 ( .a(destination_floor_elevator2[13]), .b(n1603), .out(n612) );
  inv U1052 ( .in(requested_floor[13]), .out(n546) );
  oai12 U1053 ( .b(n1603), .c(n548), .a(n613), .out(N322) );
  nand2 U1054 ( .a(destination_floor_elevator2[12]), .b(n1603), .out(n613) );
  inv U1055 ( .in(requested_floor[12]), .out(n548) );
  oai12 U1056 ( .b(n1603), .c(n555), .a(n614), .out(N321) );
  nand2 U1057 ( .a(destination_floor_elevator2[11]), .b(n1604), .out(n614) );
  inv U1058 ( .in(requested_floor[11]), .out(n555) );
  oai12 U1059 ( .b(n1604), .c(n568), .a(n615), .out(N320) );
  nand2 U1060 ( .a(destination_floor_elevator2[10]), .b(n1604), .out(n615) );
  inv U1061 ( .in(requested_floor[10]), .out(n568) );
  oai12 U1062 ( .b(n1649), .c(n616), .a(n617), .out(N32) );
  nand2 U1063 ( .a(destination_floor_elevator1[6]), .b(n1649), .out(n617) );
  oai12 U1064 ( .b(n1604), .c(n580), .a(n618), .out(N319) );
  nand2 U1065 ( .a(n1604), .b(destination_floor_elevator2[9]), .out(n618) );
  inv U1066 ( .in(requested_floor[9]), .out(n580) );
  oai12 U1067 ( .b(n1604), .c(n592), .a(n619), .out(N318) );
  nand2 U1068 ( .a(destination_floor_elevator2[8]), .b(n1604), .out(n619) );
  inv U1069 ( .in(requested_floor[8]), .out(n592) );
  oai12 U1070 ( .b(n1604), .c(n604), .a(n620), .out(N317) );
  nand2 U1071 ( .a(destination_floor_elevator2[7]), .b(n1604), .out(n620) );
  inv U1072 ( .in(requested_floor[7]), .out(n604) );
  oai12 U1073 ( .b(n1604), .c(n616), .a(n621), .out(N316) );
  nand2 U1074 ( .a(destination_floor_elevator2[6]), .b(n1604), .out(n621) );
  inv U1075 ( .in(requested_floor[6]), .out(n616) );
  oai12 U1076 ( .b(n1604), .c(n622), .a(n623), .out(N315) );
  nand2 U1077 ( .a(destination_floor_elevator2[5]), .b(n1605), .out(n623) );
  oai12 U1078 ( .b(n1605), .c(n624), .a(n625), .out(N314) );
  nand2 U1079 ( .a(destination_floor_elevator2[4]), .b(n1605), .out(n625) );
  oai12 U1080 ( .b(n1605), .c(n626), .a(n627), .out(N313) );
  nand2 U1081 ( .a(destination_floor_elevator2[3]), .b(n1605), .out(n627) );
  oai12 U1082 ( .b(n1605), .c(n628), .a(n629), .out(N312) );
  nand2 U1083 ( .a(destination_floor_elevator2[2]), .b(n1605), .out(n629) );
  oai12 U1084 ( .b(n1605), .c(n630), .a(n631), .out(N311) );
  nand2 U1085 ( .a(destination_floor_elevator2[1]), .b(n1605), .out(n631) );
  oai12 U1086 ( .b(n1605), .c(n632), .a(n633), .out(N310) );
  nand2 U1087 ( .a(destination_floor_elevator2[0]), .b(n1605), .out(n633) );
  oai12 U1088 ( .b(n1649), .c(n622), .a(n634), .out(N31) );
  nand2 U1089 ( .a(destination_floor_elevator1[5]), .b(n1650), .out(n634) );
  inv U1090 ( .in(requested_floor[5]), .out(n622) );
  oai12 U1091 ( .b(n1650), .c(n624), .a(n635), .out(N30) );
  nand2 U1092 ( .a(destination_floor_elevator1[4]), .b(n1650), .out(n635) );
  inv U1093 ( .in(requested_floor[4]), .out(n624) );
  oai12 U1094 ( .b(n1650), .c(n626), .a(n636), .out(N29) );
  nand2 U1095 ( .a(destination_floor_elevator1[3]), .b(n1650), .out(n636) );
  inv U1096 ( .in(requested_floor[3]), .out(n626) );
  oai12 U1097 ( .b(n1650), .c(n628), .a(n637), .out(N28) );
  nand2 U1098 ( .a(destination_floor_elevator1[2]), .b(n1650), .out(n637) );
  inv U1099 ( .in(requested_floor[2]), .out(n628) );
  oai12 U1100 ( .b(n1650), .c(n630), .a(n638), .out(N27) );
  nand2 U1101 ( .a(destination_floor_elevator1[1]), .b(n1650), .out(n638) );
  inv U1102 ( .in(requested_floor[1]), .out(n630) );
  oai12 U1103 ( .b(n1650), .c(n632), .a(n639), .out(N26) );
  nand2 U1104 ( .a(destination_floor_elevator1[0]), .b(n1650), .out(n639) );
  inv U1105 ( .in(requested_floor[0]), .out(n632) );
  nand2 U1106 ( .a(n775), .b(n774), .out(N154) );
  nand2 U1107 ( .a(n771), .b(n770), .out(N153) );
  nand2 U1108 ( .a(n773), .b(n772), .out(N152) );
  nand2 U1109 ( .a(n777), .b(n776), .out(N151) );
  nand2 U1110 ( .a(n779), .b(n778), .out(N150) );
  nand2 U1111 ( .a(n781), .b(n780), .out(N149) );
  nand2 U1112 ( .a(n783), .b(n782), .out(N148) );
  nand2 U1113 ( .a(n785), .b(n784), .out(N147) );
  nand2 U1114 ( .a(n787), .b(n786), .out(N146) );
  nand2 U1115 ( .a(n789), .b(n788), .out(N145) );
  nand2 U1116 ( .a(n791), .b(n790), .out(N144) );
  nand2 U1117 ( .a(n793), .b(n792), .out(N143) );
  nand2 U1118 ( .a(n795), .b(n794), .out(N142) );
  nand2 U1119 ( .a(n797), .b(n796), .out(N141) );
  nand2 U1120 ( .a(n799), .b(n798), .out(N140) );
  nand2 U1121 ( .a(n801), .b(n800), .out(N139) );
  nand2 U1122 ( .a(n803), .b(n802), .out(N138) );
  nand2 U1123 ( .a(n805), .b(n804), .out(N137) );
  nand2 U1124 ( .a(n807), .b(n806), .out(N136) );
  nand2 U1125 ( .a(n809), .b(n808), .out(N135) );
  nand2 U1126 ( .a(n811), .b(n810), .out(N134) );
  nand2 U1127 ( .a(n813), .b(n812), .out(N133) );
  nand2 U1128 ( .a(n815), .b(n814), .out(N132) );
  nand2 U1129 ( .a(n817), .b(n816), .out(N131) );
  nand2 U1130 ( .a(n819), .b(n818), .out(N130) );
  nand2 U1131 ( .a(n821), .b(n820), .out(N129) );
  nand2 U1132 ( .a(n823), .b(n822), .out(N128) );
  nand2 U1133 ( .a(n825), .b(n824), .out(N127) );
  nand2 U1134 ( .a(n827), .b(n826), .out(N126) );
  nand2 U1135 ( .a(n829), .b(n828), .out(N125) );
  nand2 U1136 ( .a(n831), .b(n830), .out(N124) );
  nand2 U1137 ( .a(n833), .b(n832), .out(N123) );
  nand2 U1138 ( .a(n835), .b(n834), .out(N122) );
  nand2 U1139 ( .a(n837), .b(n836), .out(N121) );
  nand2 U1140 ( .a(n839), .b(n838), .out(N120) );
  nand2 U1141 ( .a(n841), .b(n840), .out(N119) );
  nand2 U1142 ( .a(n843), .b(n842), .out(N118) );
  nand2 U1143 ( .a(n845), .b(n844), .out(N117) );
  nand2 U1144 ( .a(n847), .b(n846), .out(N116) );
  nand2 U1145 ( .a(n849), .b(n848), .out(N115) );
  nand2 U1146 ( .a(n851), .b(n850), .out(N114) );
  nand2 U1147 ( .a(n853), .b(n852), .out(N113) );
  nand2 U1148 ( .a(n855), .b(n854), .out(N112) );
  nand2 U1149 ( .a(n857), .b(n856), .out(N111) );
  nand2 U1150 ( .a(n859), .b(n858), .out(N110) );
  nand2 U1151 ( .a(n861), .b(n860), .out(N109) );
  nand2 U1152 ( .a(n863), .b(n862), .out(N108) );
  nand2 U1153 ( .a(n865), .b(n864), .out(N107) );
  nand2 U1154 ( .a(n867), .b(n866), .out(N106) );
  nand2 U1155 ( .a(n869), .b(n868), .out(N105) );
  nand2 U1156 ( .a(n871), .b(n870), .out(N104) );
  nand2 U1157 ( .a(n873), .b(n872), .out(N103) );
  nand2 U1158 ( .a(n875), .b(n874), .out(N102) );
  nand2 U1159 ( .a(n877), .b(n876), .out(N101) );
  nand2 U1160 ( .a(n879), .b(n878), .out(N100) );
  nor2 U1163 ( .a(n1170), .b(n1169), .out(N514) );
  nand2 U1164 ( .a(n1167), .b(n1168), .out(n1170) );
  nor2 U1165 ( .a(n1172), .b(n1171), .out(N230) );
  nand2 U1166 ( .a(n1165), .b(n1166), .out(n1172) );
  inv U1167 ( .in(n1173), .out(N607) );
  inv U1168 ( .in(n1174), .out(N609) );
  nor2 \r126/UEQ  ( .a(N505), .b(N507), .out(N509) );
  nand2 \r126/UNGT0  ( .a(N502), .b(n2842), .out(n2841) );
  nand2 \r126/UNLT0  ( .a(N438), .b(n2840), .out(n2839) );
  xor2 \r126/UEQI  ( .a(\r126/SA ), .b(\r126/SB ), .out(n2838) );
  nand2 \r126/UGTI0  ( .a(n2837), .b(\r126/SA ), .out(\r126/GTV1 [63]) );
  nand2 \r126/UGTI1  ( .a(\r126/AEQB [63]), .b(\r126/GTV [63]), .out(
        \r126/GTV2 [63]) );
  nand2 \r126/UGTI2  ( .a(\r126/GTV1 [63]), .b(\r126/GTV2 [63]), .out(N505) );
  nand2 \r126/ULTI0  ( .a(n2836), .b(\r126/SB ), .out(\r126/LTV1 [63]) );
  nand2 \r126/ULTI1  ( .a(\r126/AEQB [63]), .b(\r126/LTV [63]), .out(
        \r126/LTV2 [63]) );
  nand2 \r126/ULTI2  ( .a(\r126/LTV1 [63]), .b(\r126/LTV2 [63]), .out(N507) );
  xor2 \r126/UEQI_1  ( .a(N501), .b(N437), .out(n2835) );
  nand2 \r126/UGTI0_1  ( .a(n2834), .b(N501), .out(\r126/GTV1 [1]) );
  nand2 \r126/UGTI1_1  ( .a(\r126/AEQB [1]), .b(\r126/GTV [1]), .out(
        \r126/GTV2 [1]) );
  nand2 \r126/UGTI2_1  ( .a(\r126/GTV1 [1]), .b(\r126/GTV2 [1]), .out(
        \r126/GTV [2]) );
  nand2 \r126/ULTI0_1  ( .a(n2833), .b(N437), .out(\r126/LTV1 [1]) );
  nand2 \r126/ULTI1_1  ( .a(\r126/AEQB [1]), .b(\r126/LTV [1]), .out(
        \r126/LTV2 [1]) );
  nand2 \r126/ULTI2_1  ( .a(\r126/LTV1 [1]), .b(\r126/LTV2 [1]), .out(
        \r126/LTV [2]) );
  xor2 \r126/UEQI_2  ( .a(N500), .b(N436), .out(n2832) );
  nand2 \r126/UGTI0_2  ( .a(n2831), .b(N500), .out(\r126/GTV1 [2]) );
  nand2 \r126/UGTI1_2  ( .a(\r126/AEQB [2]), .b(\r126/GTV [2]), .out(
        \r126/GTV2 [2]) );
  nand2 \r126/UGTI2_2  ( .a(\r126/GTV1 [2]), .b(\r126/GTV2 [2]), .out(
        \r126/GTV [3]) );
  nand2 \r126/ULTI0_2  ( .a(n2830), .b(N436), .out(\r126/LTV1 [2]) );
  nand2 \r126/ULTI1_2  ( .a(\r126/AEQB [2]), .b(\r126/LTV [2]), .out(
        \r126/LTV2 [2]) );
  nand2 \r126/ULTI2_2  ( .a(\r126/LTV1 [2]), .b(\r126/LTV2 [2]), .out(
        \r126/LTV [3]) );
  xor2 \r126/UEQI_3  ( .a(N499), .b(N435), .out(n2829) );
  nand2 \r126/UGTI0_3  ( .a(n2828), .b(N499), .out(\r126/GTV1 [3]) );
  nand2 \r126/UGTI1_3  ( .a(\r126/AEQB [3]), .b(\r126/GTV [3]), .out(
        \r126/GTV2 [3]) );
  nand2 \r126/UGTI2_3  ( .a(\r126/GTV1 [3]), .b(\r126/GTV2 [3]), .out(
        \r126/GTV [4]) );
  nand2 \r126/ULTI0_3  ( .a(n2827), .b(N435), .out(\r126/LTV1 [3]) );
  nand2 \r126/ULTI1_3  ( .a(\r126/AEQB [3]), .b(\r126/LTV [3]), .out(
        \r126/LTV2 [3]) );
  nand2 \r126/ULTI2_3  ( .a(\r126/LTV1 [3]), .b(\r126/LTV2 [3]), .out(
        \r126/LTV [4]) );
  xor2 \r126/UEQI_4  ( .a(N498), .b(N434), .out(n2826) );
  nand2 \r126/UGTI0_4  ( .a(n2825), .b(N498), .out(\r126/GTV1 [4]) );
  nand2 \r126/UGTI1_4  ( .a(\r126/AEQB [4]), .b(\r126/GTV [4]), .out(
        \r126/GTV2 [4]) );
  nand2 \r126/UGTI2_4  ( .a(\r126/GTV1 [4]), .b(\r126/GTV2 [4]), .out(
        \r126/GTV [5]) );
  nand2 \r126/ULTI0_4  ( .a(n2824), .b(N434), .out(\r126/LTV1 [4]) );
  nand2 \r126/ULTI1_4  ( .a(\r126/AEQB [4]), .b(\r126/LTV [4]), .out(
        \r126/LTV2 [4]) );
  nand2 \r126/ULTI2_4  ( .a(\r126/LTV1 [4]), .b(\r126/LTV2 [4]), .out(
        \r126/LTV [5]) );
  xor2 \r126/UEQI_5  ( .a(N497), .b(N433), .out(n2823) );
  nand2 \r126/UGTI0_5  ( .a(n2822), .b(N497), .out(\r126/GTV1 [5]) );
  nand2 \r126/UGTI1_5  ( .a(\r126/AEQB [5]), .b(\r126/GTV [5]), .out(
        \r126/GTV2 [5]) );
  nand2 \r126/UGTI2_5  ( .a(\r126/GTV1 [5]), .b(\r126/GTV2 [5]), .out(
        \r126/GTV [6]) );
  nand2 \r126/ULTI0_5  ( .a(n2821), .b(N433), .out(\r126/LTV1 [5]) );
  nand2 \r126/ULTI1_5  ( .a(\r126/AEQB [5]), .b(\r126/LTV [5]), .out(
        \r126/LTV2 [5]) );
  nand2 \r126/ULTI2_5  ( .a(\r126/LTV1 [5]), .b(\r126/LTV2 [5]), .out(
        \r126/LTV [6]) );
  xor2 \r126/UEQI_6  ( .a(N496), .b(N432), .out(n2820) );
  nand2 \r126/UGTI0_6  ( .a(n2819), .b(N496), .out(\r126/GTV1 [6]) );
  nand2 \r126/UGTI1_6  ( .a(\r126/AEQB [6]), .b(\r126/GTV [6]), .out(
        \r126/GTV2 [6]) );
  nand2 \r126/UGTI2_6  ( .a(\r126/GTV1 [6]), .b(\r126/GTV2 [6]), .out(
        \r126/GTV [7]) );
  nand2 \r126/ULTI0_6  ( .a(n2818), .b(N432), .out(\r126/LTV1 [6]) );
  nand2 \r126/ULTI1_6  ( .a(\r126/AEQB [6]), .b(\r126/LTV [6]), .out(
        \r126/LTV2 [6]) );
  nand2 \r126/ULTI2_6  ( .a(\r126/LTV1 [6]), .b(\r126/LTV2 [6]), .out(
        \r126/LTV [7]) );
  xor2 \r126/UEQI_7  ( .a(N495), .b(N431), .out(n2817) );
  nand2 \r126/UGTI0_7  ( .a(n2816), .b(N495), .out(\r126/GTV1 [7]) );
  nand2 \r126/UGTI1_7  ( .a(\r126/AEQB [7]), .b(\r126/GTV [7]), .out(
        \r126/GTV2 [7]) );
  nand2 \r126/UGTI2_7  ( .a(\r126/GTV1 [7]), .b(\r126/GTV2 [7]), .out(
        \r126/GTV [8]) );
  nand2 \r126/ULTI0_7  ( .a(n2815), .b(N431), .out(\r126/LTV1 [7]) );
  nand2 \r126/ULTI1_7  ( .a(\r126/AEQB [7]), .b(\r126/LTV [7]), .out(
        \r126/LTV2 [7]) );
  nand2 \r126/ULTI2_7  ( .a(\r126/LTV1 [7]), .b(\r126/LTV2 [7]), .out(
        \r126/LTV [8]) );
  xor2 \r126/UEQI_8  ( .a(N494), .b(N430), .out(n2814) );
  nand2 \r126/UGTI0_8  ( .a(n2813), .b(N494), .out(\r126/GTV1 [8]) );
  nand2 \r126/UGTI1_8  ( .a(\r126/AEQB [8]), .b(\r126/GTV [8]), .out(
        \r126/GTV2 [8]) );
  nand2 \r126/UGTI2_8  ( .a(\r126/GTV1 [8]), .b(\r126/GTV2 [8]), .out(
        \r126/GTV [9]) );
  nand2 \r126/ULTI0_8  ( .a(n2812), .b(N430), .out(\r126/LTV1 [8]) );
  nand2 \r126/ULTI1_8  ( .a(\r126/AEQB [8]), .b(\r126/LTV [8]), .out(
        \r126/LTV2 [8]) );
  nand2 \r126/ULTI2_8  ( .a(\r126/LTV1 [8]), .b(\r126/LTV2 [8]), .out(
        \r126/LTV [9]) );
  xor2 \r126/UEQI_9  ( .a(N493), .b(N429), .out(n2811) );
  nand2 \r126/UGTI0_9  ( .a(n2810), .b(N493), .out(\r126/GTV1 [9]) );
  nand2 \r126/UGTI1_9  ( .a(\r126/AEQB [9]), .b(\r126/GTV [9]), .out(
        \r126/GTV2 [9]) );
  nand2 \r126/UGTI2_9  ( .a(\r126/GTV1 [9]), .b(\r126/GTV2 [9]), .out(
        \r126/GTV [10]) );
  nand2 \r126/ULTI0_9  ( .a(n2809), .b(N429), .out(\r126/LTV1 [9]) );
  nand2 \r126/ULTI1_9  ( .a(\r126/AEQB [9]), .b(\r126/LTV [9]), .out(
        \r126/LTV2 [9]) );
  nand2 \r126/ULTI2_9  ( .a(\r126/LTV1 [9]), .b(\r126/LTV2 [9]), .out(
        \r126/LTV [10]) );
  xor2 \r126/UEQI_10  ( .a(N492), .b(N428), .out(n2808) );
  nand2 \r126/UGTI0_10  ( .a(n2807), .b(N492), .out(\r126/GTV1 [10]) );
  nand2 \r126/UGTI1_10  ( .a(\r126/AEQB [10]), .b(\r126/GTV [10]), .out(
        \r126/GTV2 [10]) );
  nand2 \r126/UGTI2_10  ( .a(\r126/GTV1 [10]), .b(\r126/GTV2 [10]), .out(
        \r126/GTV [11]) );
  nand2 \r126/ULTI0_10  ( .a(n2806), .b(N428), .out(\r126/LTV1 [10]) );
  nand2 \r126/ULTI1_10  ( .a(\r126/AEQB [10]), .b(\r126/LTV [10]), .out(
        \r126/LTV2 [10]) );
  nand2 \r126/ULTI2_10  ( .a(\r126/LTV1 [10]), .b(\r126/LTV2 [10]), .out(
        \r126/LTV [11]) );
  xor2 \r126/UEQI_11  ( .a(N491), .b(N427), .out(n2805) );
  nand2 \r126/UGTI0_11  ( .a(n2804), .b(N491), .out(\r126/GTV1 [11]) );
  nand2 \r126/UGTI1_11  ( .a(\r126/AEQB [11]), .b(\r126/GTV [11]), .out(
        \r126/GTV2 [11]) );
  nand2 \r126/UGTI2_11  ( .a(\r126/GTV1 [11]), .b(\r126/GTV2 [11]), .out(
        \r126/GTV [12]) );
  nand2 \r126/ULTI0_11  ( .a(n2803), .b(N427), .out(\r126/LTV1 [11]) );
  nand2 \r126/ULTI1_11  ( .a(\r126/AEQB [11]), .b(\r126/LTV [11]), .out(
        \r126/LTV2 [11]) );
  nand2 \r126/ULTI2_11  ( .a(\r126/LTV1 [11]), .b(\r126/LTV2 [11]), .out(
        \r126/LTV [12]) );
  xor2 \r126/UEQI_12  ( .a(N490), .b(N426), .out(n2802) );
  nand2 \r126/UGTI0_12  ( .a(n2801), .b(N490), .out(\r126/GTV1 [12]) );
  nand2 \r126/UGTI1_12  ( .a(\r126/AEQB [12]), .b(\r126/GTV [12]), .out(
        \r126/GTV2 [12]) );
  nand2 \r126/UGTI2_12  ( .a(\r126/GTV1 [12]), .b(\r126/GTV2 [12]), .out(
        \r126/GTV [13]) );
  nand2 \r126/ULTI0_12  ( .a(n2800), .b(N426), .out(\r126/LTV1 [12]) );
  nand2 \r126/ULTI1_12  ( .a(\r126/AEQB [12]), .b(\r126/LTV [12]), .out(
        \r126/LTV2 [12]) );
  nand2 \r126/ULTI2_12  ( .a(\r126/LTV1 [12]), .b(\r126/LTV2 [12]), .out(
        \r126/LTV [13]) );
  xor2 \r126/UEQI_13  ( .a(N489), .b(N425), .out(n2799) );
  nand2 \r126/UGTI0_13  ( .a(n2798), .b(N489), .out(\r126/GTV1 [13]) );
  nand2 \r126/UGTI1_13  ( .a(\r126/AEQB [13]), .b(\r126/GTV [13]), .out(
        \r126/GTV2 [13]) );
  nand2 \r126/UGTI2_13  ( .a(\r126/GTV1 [13]), .b(\r126/GTV2 [13]), .out(
        \r126/GTV [14]) );
  nand2 \r126/ULTI0_13  ( .a(n2797), .b(N425), .out(\r126/LTV1 [13]) );
  nand2 \r126/ULTI1_13  ( .a(\r126/AEQB [13]), .b(\r126/LTV [13]), .out(
        \r126/LTV2 [13]) );
  nand2 \r126/ULTI2_13  ( .a(\r126/LTV1 [13]), .b(\r126/LTV2 [13]), .out(
        \r126/LTV [14]) );
  xor2 \r126/UEQI_14  ( .a(N488), .b(N424), .out(n2796) );
  nand2 \r126/UGTI0_14  ( .a(n2795), .b(N488), .out(\r126/GTV1 [14]) );
  nand2 \r126/UGTI1_14  ( .a(\r126/AEQB [14]), .b(\r126/GTV [14]), .out(
        \r126/GTV2 [14]) );
  nand2 \r126/UGTI2_14  ( .a(\r126/GTV1 [14]), .b(\r126/GTV2 [14]), .out(
        \r126/GTV [15]) );
  nand2 \r126/ULTI0_14  ( .a(n2794), .b(N424), .out(\r126/LTV1 [14]) );
  nand2 \r126/ULTI1_14  ( .a(\r126/AEQB [14]), .b(\r126/LTV [14]), .out(
        \r126/LTV2 [14]) );
  nand2 \r126/ULTI2_14  ( .a(\r126/LTV1 [14]), .b(\r126/LTV2 [14]), .out(
        \r126/LTV [15]) );
  xor2 \r126/UEQI_15  ( .a(N487), .b(N423), .out(n2793) );
  nand2 \r126/UGTI0_15  ( .a(n2792), .b(N487), .out(\r126/GTV1 [15]) );
  nand2 \r126/UGTI1_15  ( .a(\r126/AEQB [15]), .b(\r126/GTV [15]), .out(
        \r126/GTV2 [15]) );
  nand2 \r126/UGTI2_15  ( .a(\r126/GTV1 [15]), .b(\r126/GTV2 [15]), .out(
        \r126/GTV [16]) );
  nand2 \r126/ULTI0_15  ( .a(n2791), .b(N423), .out(\r126/LTV1 [15]) );
  nand2 \r126/ULTI1_15  ( .a(\r126/AEQB [15]), .b(\r126/LTV [15]), .out(
        \r126/LTV2 [15]) );
  nand2 \r126/ULTI2_15  ( .a(\r126/LTV1 [15]), .b(\r126/LTV2 [15]), .out(
        \r126/LTV [16]) );
  xor2 \r126/UEQI_16  ( .a(N486), .b(N422), .out(n2790) );
  nand2 \r126/UGTI0_16  ( .a(n2789), .b(N486), .out(\r126/GTV1 [16]) );
  nand2 \r126/UGTI1_16  ( .a(\r126/AEQB [16]), .b(\r126/GTV [16]), .out(
        \r126/GTV2 [16]) );
  nand2 \r126/UGTI2_16  ( .a(\r126/GTV1 [16]), .b(\r126/GTV2 [16]), .out(
        \r126/GTV [17]) );
  nand2 \r126/ULTI0_16  ( .a(n2788), .b(N422), .out(\r126/LTV1 [16]) );
  nand2 \r126/ULTI1_16  ( .a(\r126/AEQB [16]), .b(\r126/LTV [16]), .out(
        \r126/LTV2 [16]) );
  nand2 \r126/ULTI2_16  ( .a(\r126/LTV1 [16]), .b(\r126/LTV2 [16]), .out(
        \r126/LTV [17]) );
  xor2 \r126/UEQI_17  ( .a(N485), .b(N421), .out(n2787) );
  nand2 \r126/UGTI0_17  ( .a(n2786), .b(N485), .out(\r126/GTV1 [17]) );
  nand2 \r126/UGTI1_17  ( .a(\r126/AEQB [17]), .b(\r126/GTV [17]), .out(
        \r126/GTV2 [17]) );
  nand2 \r126/UGTI2_17  ( .a(\r126/GTV1 [17]), .b(\r126/GTV2 [17]), .out(
        \r126/GTV [18]) );
  nand2 \r126/ULTI0_17  ( .a(n2785), .b(N421), .out(\r126/LTV1 [17]) );
  nand2 \r126/ULTI1_17  ( .a(\r126/AEQB [17]), .b(\r126/LTV [17]), .out(
        \r126/LTV2 [17]) );
  nand2 \r126/ULTI2_17  ( .a(\r126/LTV1 [17]), .b(\r126/LTV2 [17]), .out(
        \r126/LTV [18]) );
  xor2 \r126/UEQI_18  ( .a(N484), .b(N420), .out(n2784) );
  nand2 \r126/UGTI0_18  ( .a(n2783), .b(N484), .out(\r126/GTV1 [18]) );
  nand2 \r126/UGTI1_18  ( .a(\r126/AEQB [18]), .b(\r126/GTV [18]), .out(
        \r126/GTV2 [18]) );
  nand2 \r126/UGTI2_18  ( .a(\r126/GTV1 [18]), .b(\r126/GTV2 [18]), .out(
        \r126/GTV [19]) );
  nand2 \r126/ULTI0_18  ( .a(n2782), .b(N420), .out(\r126/LTV1 [18]) );
  nand2 \r126/ULTI1_18  ( .a(\r126/AEQB [18]), .b(\r126/LTV [18]), .out(
        \r126/LTV2 [18]) );
  nand2 \r126/ULTI2_18  ( .a(\r126/LTV1 [18]), .b(\r126/LTV2 [18]), .out(
        \r126/LTV [19]) );
  xor2 \r126/UEQI_19  ( .a(N483), .b(N419), .out(n2781) );
  nand2 \r126/UGTI0_19  ( .a(n2780), .b(N483), .out(\r126/GTV1 [19]) );
  nand2 \r126/UGTI1_19  ( .a(\r126/AEQB [19]), .b(\r126/GTV [19]), .out(
        \r126/GTV2 [19]) );
  nand2 \r126/UGTI2_19  ( .a(\r126/GTV1 [19]), .b(\r126/GTV2 [19]), .out(
        \r126/GTV [20]) );
  nand2 \r126/ULTI0_19  ( .a(n2779), .b(N419), .out(\r126/LTV1 [19]) );
  nand2 \r126/ULTI1_19  ( .a(\r126/AEQB [19]), .b(\r126/LTV [19]), .out(
        \r126/LTV2 [19]) );
  nand2 \r126/ULTI2_19  ( .a(\r126/LTV1 [19]), .b(\r126/LTV2 [19]), .out(
        \r126/LTV [20]) );
  xor2 \r126/UEQI_20  ( .a(N482), .b(N418), .out(n2778) );
  nand2 \r126/UGTI0_20  ( .a(n2777), .b(N482), .out(\r126/GTV1 [20]) );
  nand2 \r126/UGTI1_20  ( .a(\r126/AEQB [20]), .b(\r126/GTV [20]), .out(
        \r126/GTV2 [20]) );
  nand2 \r126/UGTI2_20  ( .a(\r126/GTV1 [20]), .b(\r126/GTV2 [20]), .out(
        \r126/GTV [21]) );
  nand2 \r126/ULTI0_20  ( .a(n2776), .b(N418), .out(\r126/LTV1 [20]) );
  nand2 \r126/ULTI1_20  ( .a(\r126/AEQB [20]), .b(\r126/LTV [20]), .out(
        \r126/LTV2 [20]) );
  nand2 \r126/ULTI2_20  ( .a(\r126/LTV1 [20]), .b(\r126/LTV2 [20]), .out(
        \r126/LTV [21]) );
  xor2 \r126/UEQI_21  ( .a(N481), .b(N417), .out(n2775) );
  nand2 \r126/UGTI0_21  ( .a(n2774), .b(N481), .out(\r126/GTV1 [21]) );
  nand2 \r126/UGTI1_21  ( .a(\r126/AEQB [21]), .b(\r126/GTV [21]), .out(
        \r126/GTV2 [21]) );
  nand2 \r126/UGTI2_21  ( .a(\r126/GTV1 [21]), .b(\r126/GTV2 [21]), .out(
        \r126/GTV [22]) );
  nand2 \r126/ULTI0_21  ( .a(n2773), .b(N417), .out(\r126/LTV1 [21]) );
  nand2 \r126/ULTI1_21  ( .a(\r126/AEQB [21]), .b(\r126/LTV [21]), .out(
        \r126/LTV2 [21]) );
  nand2 \r126/ULTI2_21  ( .a(\r126/LTV1 [21]), .b(\r126/LTV2 [21]), .out(
        \r126/LTV [22]) );
  xor2 \r126/UEQI_22  ( .a(N480), .b(N416), .out(n2772) );
  nand2 \r126/UGTI0_22  ( .a(n2771), .b(N480), .out(\r126/GTV1 [22]) );
  nand2 \r126/UGTI1_22  ( .a(\r126/AEQB [22]), .b(\r126/GTV [22]), .out(
        \r126/GTV2 [22]) );
  nand2 \r126/UGTI2_22  ( .a(\r126/GTV1 [22]), .b(\r126/GTV2 [22]), .out(
        \r126/GTV [23]) );
  nand2 \r126/ULTI0_22  ( .a(n2770), .b(N416), .out(\r126/LTV1 [22]) );
  nand2 \r126/ULTI1_22  ( .a(\r126/AEQB [22]), .b(\r126/LTV [22]), .out(
        \r126/LTV2 [22]) );
  nand2 \r126/ULTI2_22  ( .a(\r126/LTV1 [22]), .b(\r126/LTV2 [22]), .out(
        \r126/LTV [23]) );
  xor2 \r126/UEQI_23  ( .a(N479), .b(N415), .out(n2769) );
  nand2 \r126/UGTI0_23  ( .a(n2768), .b(N479), .out(\r126/GTV1 [23]) );
  nand2 \r126/UGTI1_23  ( .a(\r126/AEQB [23]), .b(\r126/GTV [23]), .out(
        \r126/GTV2 [23]) );
  nand2 \r126/UGTI2_23  ( .a(\r126/GTV1 [23]), .b(\r126/GTV2 [23]), .out(
        \r126/GTV [24]) );
  nand2 \r126/ULTI0_23  ( .a(n2767), .b(N415), .out(\r126/LTV1 [23]) );
  nand2 \r126/ULTI1_23  ( .a(\r126/AEQB [23]), .b(\r126/LTV [23]), .out(
        \r126/LTV2 [23]) );
  nand2 \r126/ULTI2_23  ( .a(\r126/LTV1 [23]), .b(\r126/LTV2 [23]), .out(
        \r126/LTV [24]) );
  xor2 \r126/UEQI_24  ( .a(N478), .b(N414), .out(n2766) );
  nand2 \r126/UGTI0_24  ( .a(n2765), .b(N478), .out(\r126/GTV1 [24]) );
  nand2 \r126/UGTI1_24  ( .a(\r126/AEQB [24]), .b(\r126/GTV [24]), .out(
        \r126/GTV2 [24]) );
  nand2 \r126/UGTI2_24  ( .a(\r126/GTV1 [24]), .b(\r126/GTV2 [24]), .out(
        \r126/GTV [25]) );
  nand2 \r126/ULTI0_24  ( .a(n2764), .b(N414), .out(\r126/LTV1 [24]) );
  nand2 \r126/ULTI1_24  ( .a(\r126/AEQB [24]), .b(\r126/LTV [24]), .out(
        \r126/LTV2 [24]) );
  nand2 \r126/ULTI2_24  ( .a(\r126/LTV1 [24]), .b(\r126/LTV2 [24]), .out(
        \r126/LTV [25]) );
  xor2 \r126/UEQI_25  ( .a(N477), .b(N413), .out(n2763) );
  nand2 \r126/UGTI0_25  ( .a(n2762), .b(N477), .out(\r126/GTV1 [25]) );
  nand2 \r126/UGTI1_25  ( .a(\r126/AEQB [25]), .b(\r126/GTV [25]), .out(
        \r126/GTV2 [25]) );
  nand2 \r126/UGTI2_25  ( .a(\r126/GTV1 [25]), .b(\r126/GTV2 [25]), .out(
        \r126/GTV [26]) );
  nand2 \r126/ULTI0_25  ( .a(n2761), .b(N413), .out(\r126/LTV1 [25]) );
  nand2 \r126/ULTI1_25  ( .a(\r126/AEQB [25]), .b(\r126/LTV [25]), .out(
        \r126/LTV2 [25]) );
  nand2 \r126/ULTI2_25  ( .a(\r126/LTV1 [25]), .b(\r126/LTV2 [25]), .out(
        \r126/LTV [26]) );
  xor2 \r126/UEQI_26  ( .a(N476), .b(N412), .out(n2760) );
  nand2 \r126/UGTI0_26  ( .a(n2759), .b(N476), .out(\r126/GTV1 [26]) );
  nand2 \r126/UGTI1_26  ( .a(\r126/AEQB [26]), .b(\r126/GTV [26]), .out(
        \r126/GTV2 [26]) );
  nand2 \r126/UGTI2_26  ( .a(\r126/GTV1 [26]), .b(\r126/GTV2 [26]), .out(
        \r126/GTV [27]) );
  nand2 \r126/ULTI0_26  ( .a(n2758), .b(N412), .out(\r126/LTV1 [26]) );
  nand2 \r126/ULTI1_26  ( .a(\r126/AEQB [26]), .b(\r126/LTV [26]), .out(
        \r126/LTV2 [26]) );
  nand2 \r126/ULTI2_26  ( .a(\r126/LTV1 [26]), .b(\r126/LTV2 [26]), .out(
        \r126/LTV [27]) );
  xor2 \r126/UEQI_27  ( .a(N475), .b(N411), .out(n2757) );
  nand2 \r126/UGTI0_27  ( .a(n2756), .b(N475), .out(\r126/GTV1 [27]) );
  nand2 \r126/UGTI1_27  ( .a(\r126/AEQB [27]), .b(\r126/GTV [27]), .out(
        \r126/GTV2 [27]) );
  nand2 \r126/UGTI2_27  ( .a(\r126/GTV1 [27]), .b(\r126/GTV2 [27]), .out(
        \r126/GTV [28]) );
  nand2 \r126/ULTI0_27  ( .a(n2755), .b(N411), .out(\r126/LTV1 [27]) );
  nand2 \r126/ULTI1_27  ( .a(\r126/AEQB [27]), .b(\r126/LTV [27]), .out(
        \r126/LTV2 [27]) );
  nand2 \r126/ULTI2_27  ( .a(\r126/LTV1 [27]), .b(\r126/LTV2 [27]), .out(
        \r126/LTV [28]) );
  xor2 \r126/UEQI_28  ( .a(N474), .b(N410), .out(n2754) );
  nand2 \r126/UGTI0_28  ( .a(n2753), .b(N474), .out(\r126/GTV1 [28]) );
  nand2 \r126/UGTI1_28  ( .a(\r126/AEQB [28]), .b(\r126/GTV [28]), .out(
        \r126/GTV2 [28]) );
  nand2 \r126/UGTI2_28  ( .a(\r126/GTV1 [28]), .b(\r126/GTV2 [28]), .out(
        \r126/GTV [29]) );
  nand2 \r126/ULTI0_28  ( .a(n2752), .b(N410), .out(\r126/LTV1 [28]) );
  nand2 \r126/ULTI1_28  ( .a(\r126/AEQB [28]), .b(\r126/LTV [28]), .out(
        \r126/LTV2 [28]) );
  nand2 \r126/ULTI2_28  ( .a(\r126/LTV1 [28]), .b(\r126/LTV2 [28]), .out(
        \r126/LTV [29]) );
  xor2 \r126/UEQI_29  ( .a(N473), .b(N409), .out(n2751) );
  nand2 \r126/UGTI0_29  ( .a(n2750), .b(N473), .out(\r126/GTV1 [29]) );
  nand2 \r126/UGTI1_29  ( .a(\r126/AEQB [29]), .b(\r126/GTV [29]), .out(
        \r126/GTV2 [29]) );
  nand2 \r126/UGTI2_29  ( .a(\r126/GTV1 [29]), .b(\r126/GTV2 [29]), .out(
        \r126/GTV [30]) );
  nand2 \r126/ULTI0_29  ( .a(n2749), .b(N409), .out(\r126/LTV1 [29]) );
  nand2 \r126/ULTI1_29  ( .a(\r126/AEQB [29]), .b(\r126/LTV [29]), .out(
        \r126/LTV2 [29]) );
  nand2 \r126/ULTI2_29  ( .a(\r126/LTV1 [29]), .b(\r126/LTV2 [29]), .out(
        \r126/LTV [30]) );
  xor2 \r126/UEQI_30  ( .a(N472), .b(N408), .out(n2748) );
  nand2 \r126/UGTI0_30  ( .a(n2747), .b(N472), .out(\r126/GTV1 [30]) );
  nand2 \r126/UGTI1_30  ( .a(\r126/AEQB [30]), .b(\r126/GTV [30]), .out(
        \r126/GTV2 [30]) );
  nand2 \r126/UGTI2_30  ( .a(\r126/GTV1 [30]), .b(\r126/GTV2 [30]), .out(
        \r126/GTV [31]) );
  nand2 \r126/ULTI0_30  ( .a(n2746), .b(N408), .out(\r126/LTV1 [30]) );
  nand2 \r126/ULTI1_30  ( .a(\r126/AEQB [30]), .b(\r126/LTV [30]), .out(
        \r126/LTV2 [30]) );
  nand2 \r126/ULTI2_30  ( .a(\r126/LTV1 [30]), .b(\r126/LTV2 [30]), .out(
        \r126/LTV [31]) );
  xor2 \r126/UEQI_31  ( .a(N471), .b(N407), .out(n2745) );
  nand2 \r126/UGTI0_31  ( .a(n2744), .b(N471), .out(\r126/GTV1 [31]) );
  nand2 \r126/UGTI1_31  ( .a(\r126/AEQB [31]), .b(\r126/GTV [31]), .out(
        \r126/GTV2 [31]) );
  nand2 \r126/UGTI2_31  ( .a(\r126/GTV1 [31]), .b(\r126/GTV2 [31]), .out(
        \r126/GTV [32]) );
  nand2 \r126/ULTI0_31  ( .a(n2743), .b(N407), .out(\r126/LTV1 [31]) );
  nand2 \r126/ULTI1_31  ( .a(\r126/AEQB [31]), .b(\r126/LTV [31]), .out(
        \r126/LTV2 [31]) );
  nand2 \r126/ULTI2_31  ( .a(\r126/LTV1 [31]), .b(\r126/LTV2 [31]), .out(
        \r126/LTV [32]) );
  xor2 \r126/UEQI_32  ( .a(N470), .b(N406), .out(n2742) );
  nand2 \r126/UGTI0_32  ( .a(n2741), .b(N470), .out(\r126/GTV1 [32]) );
  nand2 \r126/UGTI1_32  ( .a(\r126/AEQB [32]), .b(\r126/GTV [32]), .out(
        \r126/GTV2 [32]) );
  nand2 \r126/UGTI2_32  ( .a(\r126/GTV1 [32]), .b(\r126/GTV2 [32]), .out(
        \r126/GTV [33]) );
  nand2 \r126/ULTI0_32  ( .a(n2740), .b(N406), .out(\r126/LTV1 [32]) );
  nand2 \r126/ULTI1_32  ( .a(\r126/AEQB [32]), .b(\r126/LTV [32]), .out(
        \r126/LTV2 [32]) );
  nand2 \r126/ULTI2_32  ( .a(\r126/LTV1 [32]), .b(\r126/LTV2 [32]), .out(
        \r126/LTV [33]) );
  xor2 \r126/UEQI_33  ( .a(N469), .b(N405), .out(n2739) );
  nand2 \r126/UGTI0_33  ( .a(n2738), .b(N469), .out(\r126/GTV1 [33]) );
  nand2 \r126/UGTI1_33  ( .a(\r126/AEQB [33]), .b(\r126/GTV [33]), .out(
        \r126/GTV2 [33]) );
  nand2 \r126/UGTI2_33  ( .a(\r126/GTV1 [33]), .b(\r126/GTV2 [33]), .out(
        \r126/GTV [34]) );
  nand2 \r126/ULTI0_33  ( .a(n2737), .b(N405), .out(\r126/LTV1 [33]) );
  nand2 \r126/ULTI1_33  ( .a(\r126/AEQB [33]), .b(\r126/LTV [33]), .out(
        \r126/LTV2 [33]) );
  nand2 \r126/ULTI2_33  ( .a(\r126/LTV1 [33]), .b(\r126/LTV2 [33]), .out(
        \r126/LTV [34]) );
  xor2 \r126/UEQI_34  ( .a(N468), .b(N404), .out(n2736) );
  nand2 \r126/UGTI0_34  ( .a(n2735), .b(N468), .out(\r126/GTV1 [34]) );
  nand2 \r126/UGTI1_34  ( .a(\r126/AEQB [34]), .b(\r126/GTV [34]), .out(
        \r126/GTV2 [34]) );
  nand2 \r126/UGTI2_34  ( .a(\r126/GTV1 [34]), .b(\r126/GTV2 [34]), .out(
        \r126/GTV [35]) );
  nand2 \r126/ULTI0_34  ( .a(n2734), .b(N404), .out(\r126/LTV1 [34]) );
  nand2 \r126/ULTI1_34  ( .a(\r126/AEQB [34]), .b(\r126/LTV [34]), .out(
        \r126/LTV2 [34]) );
  nand2 \r126/ULTI2_34  ( .a(\r126/LTV1 [34]), .b(\r126/LTV2 [34]), .out(
        \r126/LTV [35]) );
  xor2 \r126/UEQI_35  ( .a(N467), .b(N403), .out(n2733) );
  nand2 \r126/UGTI0_35  ( .a(n2732), .b(N467), .out(\r126/GTV1 [35]) );
  nand2 \r126/UGTI1_35  ( .a(\r126/AEQB [35]), .b(\r126/GTV [35]), .out(
        \r126/GTV2 [35]) );
  nand2 \r126/UGTI2_35  ( .a(\r126/GTV1 [35]), .b(\r126/GTV2 [35]), .out(
        \r126/GTV [36]) );
  nand2 \r126/ULTI0_35  ( .a(n2731), .b(N403), .out(\r126/LTV1 [35]) );
  nand2 \r126/ULTI1_35  ( .a(\r126/AEQB [35]), .b(\r126/LTV [35]), .out(
        \r126/LTV2 [35]) );
  nand2 \r126/ULTI2_35  ( .a(\r126/LTV1 [35]), .b(\r126/LTV2 [35]), .out(
        \r126/LTV [36]) );
  xor2 \r126/UEQI_36  ( .a(N466), .b(N402), .out(n2730) );
  nand2 \r126/UGTI0_36  ( .a(n2729), .b(N466), .out(\r126/GTV1 [36]) );
  nand2 \r126/UGTI1_36  ( .a(\r126/AEQB [36]), .b(\r126/GTV [36]), .out(
        \r126/GTV2 [36]) );
  nand2 \r126/UGTI2_36  ( .a(\r126/GTV1 [36]), .b(\r126/GTV2 [36]), .out(
        \r126/GTV [37]) );
  nand2 \r126/ULTI0_36  ( .a(n2728), .b(N402), .out(\r126/LTV1 [36]) );
  nand2 \r126/ULTI1_36  ( .a(\r126/AEQB [36]), .b(\r126/LTV [36]), .out(
        \r126/LTV2 [36]) );
  nand2 \r126/ULTI2_36  ( .a(\r126/LTV1 [36]), .b(\r126/LTV2 [36]), .out(
        \r126/LTV [37]) );
  xor2 \r126/UEQI_37  ( .a(N465), .b(N401), .out(n2727) );
  nand2 \r126/UGTI0_37  ( .a(n2726), .b(N465), .out(\r126/GTV1 [37]) );
  nand2 \r126/UGTI1_37  ( .a(\r126/AEQB [37]), .b(\r126/GTV [37]), .out(
        \r126/GTV2 [37]) );
  nand2 \r126/UGTI2_37  ( .a(\r126/GTV1 [37]), .b(\r126/GTV2 [37]), .out(
        \r126/GTV [38]) );
  nand2 \r126/ULTI0_37  ( .a(n2725), .b(N401), .out(\r126/LTV1 [37]) );
  nand2 \r126/ULTI1_37  ( .a(\r126/AEQB [37]), .b(\r126/LTV [37]), .out(
        \r126/LTV2 [37]) );
  nand2 \r126/ULTI2_37  ( .a(\r126/LTV1 [37]), .b(\r126/LTV2 [37]), .out(
        \r126/LTV [38]) );
  xor2 \r126/UEQI_38  ( .a(N464), .b(N400), .out(n2724) );
  nand2 \r126/UGTI0_38  ( .a(n2723), .b(N464), .out(\r126/GTV1 [38]) );
  nand2 \r126/UGTI1_38  ( .a(\r126/AEQB [38]), .b(\r126/GTV [38]), .out(
        \r126/GTV2 [38]) );
  nand2 \r126/UGTI2_38  ( .a(\r126/GTV1 [38]), .b(\r126/GTV2 [38]), .out(
        \r126/GTV [39]) );
  nand2 \r126/ULTI0_38  ( .a(n2722), .b(N400), .out(\r126/LTV1 [38]) );
  nand2 \r126/ULTI1_38  ( .a(\r126/AEQB [38]), .b(\r126/LTV [38]), .out(
        \r126/LTV2 [38]) );
  nand2 \r126/ULTI2_38  ( .a(\r126/LTV1 [38]), .b(\r126/LTV2 [38]), .out(
        \r126/LTV [39]) );
  xor2 \r126/UEQI_39  ( .a(N463), .b(N399), .out(n2721) );
  nand2 \r126/UGTI0_39  ( .a(n2720), .b(N463), .out(\r126/GTV1 [39]) );
  nand2 \r126/UGTI1_39  ( .a(\r126/AEQB [39]), .b(\r126/GTV [39]), .out(
        \r126/GTV2 [39]) );
  nand2 \r126/UGTI2_39  ( .a(\r126/GTV1 [39]), .b(\r126/GTV2 [39]), .out(
        \r126/GTV [40]) );
  nand2 \r126/ULTI0_39  ( .a(n2719), .b(N399), .out(\r126/LTV1 [39]) );
  nand2 \r126/ULTI1_39  ( .a(\r126/AEQB [39]), .b(\r126/LTV [39]), .out(
        \r126/LTV2 [39]) );
  nand2 \r126/ULTI2_39  ( .a(\r126/LTV1 [39]), .b(\r126/LTV2 [39]), .out(
        \r126/LTV [40]) );
  xor2 \r126/UEQI_40  ( .a(N462), .b(N398), .out(n2718) );
  nand2 \r126/UGTI0_40  ( .a(n2717), .b(N462), .out(\r126/GTV1 [40]) );
  nand2 \r126/UGTI1_40  ( .a(\r126/AEQB [40]), .b(\r126/GTV [40]), .out(
        \r126/GTV2 [40]) );
  nand2 \r126/UGTI2_40  ( .a(\r126/GTV1 [40]), .b(\r126/GTV2 [40]), .out(
        \r126/GTV [41]) );
  nand2 \r126/ULTI0_40  ( .a(n2716), .b(N398), .out(\r126/LTV1 [40]) );
  nand2 \r126/ULTI1_40  ( .a(\r126/AEQB [40]), .b(\r126/LTV [40]), .out(
        \r126/LTV2 [40]) );
  nand2 \r126/ULTI2_40  ( .a(\r126/LTV1 [40]), .b(\r126/LTV2 [40]), .out(
        \r126/LTV [41]) );
  xor2 \r126/UEQI_41  ( .a(N461), .b(N397), .out(n2715) );
  nand2 \r126/UGTI0_41  ( .a(n2714), .b(N461), .out(\r126/GTV1 [41]) );
  nand2 \r126/UGTI1_41  ( .a(\r126/AEQB [41]), .b(\r126/GTV [41]), .out(
        \r126/GTV2 [41]) );
  nand2 \r126/UGTI2_41  ( .a(\r126/GTV1 [41]), .b(\r126/GTV2 [41]), .out(
        \r126/GTV [42]) );
  nand2 \r126/ULTI0_41  ( .a(n2713), .b(N397), .out(\r126/LTV1 [41]) );
  nand2 \r126/ULTI1_41  ( .a(\r126/AEQB [41]), .b(\r126/LTV [41]), .out(
        \r126/LTV2 [41]) );
  nand2 \r126/ULTI2_41  ( .a(\r126/LTV1 [41]), .b(\r126/LTV2 [41]), .out(
        \r126/LTV [42]) );
  xor2 \r126/UEQI_42  ( .a(N460), .b(N396), .out(n2712) );
  nand2 \r126/UGTI0_42  ( .a(n2711), .b(N460), .out(\r126/GTV1 [42]) );
  nand2 \r126/UGTI1_42  ( .a(\r126/AEQB [42]), .b(\r126/GTV [42]), .out(
        \r126/GTV2 [42]) );
  nand2 \r126/UGTI2_42  ( .a(\r126/GTV1 [42]), .b(\r126/GTV2 [42]), .out(
        \r126/GTV [43]) );
  nand2 \r126/ULTI0_42  ( .a(n2710), .b(N396), .out(\r126/LTV1 [42]) );
  nand2 \r126/ULTI1_42  ( .a(\r126/AEQB [42]), .b(\r126/LTV [42]), .out(
        \r126/LTV2 [42]) );
  nand2 \r126/ULTI2_42  ( .a(\r126/LTV1 [42]), .b(\r126/LTV2 [42]), .out(
        \r126/LTV [43]) );
  xor2 \r126/UEQI_43  ( .a(N459), .b(N395), .out(n2709) );
  nand2 \r126/UGTI0_43  ( .a(n2708), .b(N459), .out(\r126/GTV1 [43]) );
  nand2 \r126/UGTI1_43  ( .a(\r126/AEQB [43]), .b(\r126/GTV [43]), .out(
        \r126/GTV2 [43]) );
  nand2 \r126/UGTI2_43  ( .a(\r126/GTV1 [43]), .b(\r126/GTV2 [43]), .out(
        \r126/GTV [44]) );
  nand2 \r126/ULTI0_43  ( .a(n2707), .b(N395), .out(\r126/LTV1 [43]) );
  nand2 \r126/ULTI1_43  ( .a(\r126/AEQB [43]), .b(\r126/LTV [43]), .out(
        \r126/LTV2 [43]) );
  nand2 \r126/ULTI2_43  ( .a(\r126/LTV1 [43]), .b(\r126/LTV2 [43]), .out(
        \r126/LTV [44]) );
  xor2 \r126/UEQI_44  ( .a(N458), .b(N394), .out(n2706) );
  nand2 \r126/UGTI0_44  ( .a(n2705), .b(N458), .out(\r126/GTV1 [44]) );
  nand2 \r126/UGTI1_44  ( .a(\r126/AEQB [44]), .b(\r126/GTV [44]), .out(
        \r126/GTV2 [44]) );
  nand2 \r126/UGTI2_44  ( .a(\r126/GTV1 [44]), .b(\r126/GTV2 [44]), .out(
        \r126/GTV [45]) );
  nand2 \r126/ULTI0_44  ( .a(n2704), .b(N394), .out(\r126/LTV1 [44]) );
  nand2 \r126/ULTI1_44  ( .a(\r126/AEQB [44]), .b(\r126/LTV [44]), .out(
        \r126/LTV2 [44]) );
  nand2 \r126/ULTI2_44  ( .a(\r126/LTV1 [44]), .b(\r126/LTV2 [44]), .out(
        \r126/LTV [45]) );
  xor2 \r126/UEQI_45  ( .a(N457), .b(N393), .out(n2703) );
  nand2 \r126/UGTI0_45  ( .a(n2702), .b(N457), .out(\r126/GTV1 [45]) );
  nand2 \r126/UGTI1_45  ( .a(\r126/AEQB [45]), .b(\r126/GTV [45]), .out(
        \r126/GTV2 [45]) );
  nand2 \r126/UGTI2_45  ( .a(\r126/GTV1 [45]), .b(\r126/GTV2 [45]), .out(
        \r126/GTV [46]) );
  nand2 \r126/ULTI0_45  ( .a(n2701), .b(N393), .out(\r126/LTV1 [45]) );
  nand2 \r126/ULTI1_45  ( .a(\r126/AEQB [45]), .b(\r126/LTV [45]), .out(
        \r126/LTV2 [45]) );
  nand2 \r126/ULTI2_45  ( .a(\r126/LTV1 [45]), .b(\r126/LTV2 [45]), .out(
        \r126/LTV [46]) );
  xor2 \r126/UEQI_46  ( .a(N456), .b(N392), .out(n2700) );
  nand2 \r126/UGTI0_46  ( .a(n2699), .b(N456), .out(\r126/GTV1 [46]) );
  nand2 \r126/UGTI1_46  ( .a(\r126/AEQB [46]), .b(\r126/GTV [46]), .out(
        \r126/GTV2 [46]) );
  nand2 \r126/UGTI2_46  ( .a(\r126/GTV1 [46]), .b(\r126/GTV2 [46]), .out(
        \r126/GTV [47]) );
  nand2 \r126/ULTI0_46  ( .a(n2698), .b(N392), .out(\r126/LTV1 [46]) );
  nand2 \r126/ULTI1_46  ( .a(\r126/AEQB [46]), .b(\r126/LTV [46]), .out(
        \r126/LTV2 [46]) );
  nand2 \r126/ULTI2_46  ( .a(\r126/LTV1 [46]), .b(\r126/LTV2 [46]), .out(
        \r126/LTV [47]) );
  xor2 \r126/UEQI_47  ( .a(N455), .b(N391), .out(n2697) );
  nand2 \r126/UGTI0_47  ( .a(n2696), .b(N455), .out(\r126/GTV1 [47]) );
  nand2 \r126/UGTI1_47  ( .a(\r126/AEQB [47]), .b(\r126/GTV [47]), .out(
        \r126/GTV2 [47]) );
  nand2 \r126/UGTI2_47  ( .a(\r126/GTV1 [47]), .b(\r126/GTV2 [47]), .out(
        \r126/GTV [48]) );
  nand2 \r126/ULTI0_47  ( .a(n2695), .b(N391), .out(\r126/LTV1 [47]) );
  nand2 \r126/ULTI1_47  ( .a(\r126/AEQB [47]), .b(\r126/LTV [47]), .out(
        \r126/LTV2 [47]) );
  nand2 \r126/ULTI2_47  ( .a(\r126/LTV1 [47]), .b(\r126/LTV2 [47]), .out(
        \r126/LTV [48]) );
  xor2 \r126/UEQI_48  ( .a(N454), .b(N390), .out(n2694) );
  nand2 \r126/UGTI0_48  ( .a(n2693), .b(N454), .out(\r126/GTV1 [48]) );
  nand2 \r126/UGTI1_48  ( .a(\r126/AEQB [48]), .b(\r126/GTV [48]), .out(
        \r126/GTV2 [48]) );
  nand2 \r126/UGTI2_48  ( .a(\r126/GTV1 [48]), .b(\r126/GTV2 [48]), .out(
        \r126/GTV [49]) );
  nand2 \r126/ULTI0_48  ( .a(n2692), .b(N390), .out(\r126/LTV1 [48]) );
  nand2 \r126/ULTI1_48  ( .a(\r126/AEQB [48]), .b(\r126/LTV [48]), .out(
        \r126/LTV2 [48]) );
  nand2 \r126/ULTI2_48  ( .a(\r126/LTV1 [48]), .b(\r126/LTV2 [48]), .out(
        \r126/LTV [49]) );
  xor2 \r126/UEQI_49  ( .a(N453), .b(N389), .out(n2691) );
  nand2 \r126/UGTI0_49  ( .a(n2690), .b(N453), .out(\r126/GTV1 [49]) );
  nand2 \r126/UGTI1_49  ( .a(\r126/AEQB [49]), .b(\r126/GTV [49]), .out(
        \r126/GTV2 [49]) );
  nand2 \r126/UGTI2_49  ( .a(\r126/GTV1 [49]), .b(\r126/GTV2 [49]), .out(
        \r126/GTV [50]) );
  nand2 \r126/ULTI0_49  ( .a(n2689), .b(N389), .out(\r126/LTV1 [49]) );
  nand2 \r126/ULTI1_49  ( .a(\r126/AEQB [49]), .b(\r126/LTV [49]), .out(
        \r126/LTV2 [49]) );
  nand2 \r126/ULTI2_49  ( .a(\r126/LTV1 [49]), .b(\r126/LTV2 [49]), .out(
        \r126/LTV [50]) );
  xor2 \r126/UEQI_50  ( .a(N452), .b(N388), .out(n2688) );
  nand2 \r126/UGTI0_50  ( .a(n2687), .b(N452), .out(\r126/GTV1 [50]) );
  nand2 \r126/UGTI1_50  ( .a(\r126/AEQB [50]), .b(\r126/GTV [50]), .out(
        \r126/GTV2 [50]) );
  nand2 \r126/UGTI2_50  ( .a(\r126/GTV1 [50]), .b(\r126/GTV2 [50]), .out(
        \r126/GTV [51]) );
  nand2 \r126/ULTI0_50  ( .a(n2686), .b(N388), .out(\r126/LTV1 [50]) );
  nand2 \r126/ULTI1_50  ( .a(\r126/AEQB [50]), .b(\r126/LTV [50]), .out(
        \r126/LTV2 [50]) );
  nand2 \r126/ULTI2_50  ( .a(\r126/LTV1 [50]), .b(\r126/LTV2 [50]), .out(
        \r126/LTV [51]) );
  xor2 \r126/UEQI_51  ( .a(N451), .b(N387), .out(n2685) );
  nand2 \r126/UGTI0_51  ( .a(n2684), .b(N451), .out(\r126/GTV1 [51]) );
  nand2 \r126/UGTI1_51  ( .a(\r126/AEQB [51]), .b(\r126/GTV [51]), .out(
        \r126/GTV2 [51]) );
  nand2 \r126/UGTI2_51  ( .a(\r126/GTV1 [51]), .b(\r126/GTV2 [51]), .out(
        \r126/GTV [52]) );
  nand2 \r126/ULTI0_51  ( .a(n2683), .b(N387), .out(\r126/LTV1 [51]) );
  nand2 \r126/ULTI1_51  ( .a(\r126/AEQB [51]), .b(\r126/LTV [51]), .out(
        \r126/LTV2 [51]) );
  nand2 \r126/ULTI2_51  ( .a(\r126/LTV1 [51]), .b(\r126/LTV2 [51]), .out(
        \r126/LTV [52]) );
  xor2 \r126/UEQI_52  ( .a(N450), .b(N386), .out(n2682) );
  nand2 \r126/UGTI0_52  ( .a(n2681), .b(N450), .out(\r126/GTV1 [52]) );
  nand2 \r126/UGTI1_52  ( .a(\r126/AEQB [52]), .b(\r126/GTV [52]), .out(
        \r126/GTV2 [52]) );
  nand2 \r126/UGTI2_52  ( .a(\r126/GTV1 [52]), .b(\r126/GTV2 [52]), .out(
        \r126/GTV [53]) );
  nand2 \r126/ULTI0_52  ( .a(n2680), .b(N386), .out(\r126/LTV1 [52]) );
  nand2 \r126/ULTI1_52  ( .a(\r126/AEQB [52]), .b(\r126/LTV [52]), .out(
        \r126/LTV2 [52]) );
  nand2 \r126/ULTI2_52  ( .a(\r126/LTV1 [52]), .b(\r126/LTV2 [52]), .out(
        \r126/LTV [53]) );
  xor2 \r126/UEQI_53  ( .a(N449), .b(N385), .out(n2679) );
  nand2 \r126/UGTI0_53  ( .a(n2678), .b(N449), .out(\r126/GTV1 [53]) );
  nand2 \r126/UGTI1_53  ( .a(\r126/AEQB [53]), .b(\r126/GTV [53]), .out(
        \r126/GTV2 [53]) );
  nand2 \r126/UGTI2_53  ( .a(\r126/GTV1 [53]), .b(\r126/GTV2 [53]), .out(
        \r126/GTV [54]) );
  nand2 \r126/ULTI0_53  ( .a(n2677), .b(N385), .out(\r126/LTV1 [53]) );
  nand2 \r126/ULTI1_53  ( .a(\r126/AEQB [53]), .b(\r126/LTV [53]), .out(
        \r126/LTV2 [53]) );
  nand2 \r126/ULTI2_53  ( .a(\r126/LTV1 [53]), .b(\r126/LTV2 [53]), .out(
        \r126/LTV [54]) );
  xor2 \r126/UEQI_54  ( .a(N448), .b(N384), .out(n2676) );
  nand2 \r126/UGTI0_54  ( .a(n2675), .b(N448), .out(\r126/GTV1 [54]) );
  nand2 \r126/UGTI1_54  ( .a(\r126/AEQB [54]), .b(\r126/GTV [54]), .out(
        \r126/GTV2 [54]) );
  nand2 \r126/UGTI2_54  ( .a(\r126/GTV1 [54]), .b(\r126/GTV2 [54]), .out(
        \r126/GTV [55]) );
  nand2 \r126/ULTI0_54  ( .a(n2674), .b(N384), .out(\r126/LTV1 [54]) );
  nand2 \r126/ULTI1_54  ( .a(\r126/AEQB [54]), .b(\r126/LTV [54]), .out(
        \r126/LTV2 [54]) );
  nand2 \r126/ULTI2_54  ( .a(\r126/LTV1 [54]), .b(\r126/LTV2 [54]), .out(
        \r126/LTV [55]) );
  xor2 \r126/UEQI_55  ( .a(N447), .b(N383), .out(n2673) );
  nand2 \r126/UGTI0_55  ( .a(n2672), .b(N447), .out(\r126/GTV1 [55]) );
  nand2 \r126/UGTI1_55  ( .a(\r126/AEQB [55]), .b(\r126/GTV [55]), .out(
        \r126/GTV2 [55]) );
  nand2 \r126/UGTI2_55  ( .a(\r126/GTV1 [55]), .b(\r126/GTV2 [55]), .out(
        \r126/GTV [56]) );
  nand2 \r126/ULTI0_55  ( .a(n2671), .b(N383), .out(\r126/LTV1 [55]) );
  nand2 \r126/ULTI1_55  ( .a(\r126/AEQB [55]), .b(\r126/LTV [55]), .out(
        \r126/LTV2 [55]) );
  nand2 \r126/ULTI2_55  ( .a(\r126/LTV1 [55]), .b(\r126/LTV2 [55]), .out(
        \r126/LTV [56]) );
  xor2 \r126/UEQI_56  ( .a(N446), .b(N382), .out(n2670) );
  nand2 \r126/UGTI0_56  ( .a(n2669), .b(N446), .out(\r126/GTV1 [56]) );
  nand2 \r126/UGTI1_56  ( .a(\r126/AEQB [56]), .b(\r126/GTV [56]), .out(
        \r126/GTV2 [56]) );
  nand2 \r126/UGTI2_56  ( .a(\r126/GTV1 [56]), .b(\r126/GTV2 [56]), .out(
        \r126/GTV [57]) );
  nand2 \r126/ULTI0_56  ( .a(n2668), .b(N382), .out(\r126/LTV1 [56]) );
  nand2 \r126/ULTI1_56  ( .a(\r126/AEQB [56]), .b(\r126/LTV [56]), .out(
        \r126/LTV2 [56]) );
  nand2 \r126/ULTI2_56  ( .a(\r126/LTV1 [56]), .b(\r126/LTV2 [56]), .out(
        \r126/LTV [57]) );
  xor2 \r126/UEQI_57  ( .a(N445), .b(N381), .out(n2667) );
  nand2 \r126/UGTI0_57  ( .a(n2666), .b(N445), .out(\r126/GTV1 [57]) );
  nand2 \r126/UGTI1_57  ( .a(\r126/AEQB [57]), .b(\r126/GTV [57]), .out(
        \r126/GTV2 [57]) );
  nand2 \r126/UGTI2_57  ( .a(\r126/GTV1 [57]), .b(\r126/GTV2 [57]), .out(
        \r126/GTV [58]) );
  nand2 \r126/ULTI0_57  ( .a(n2665), .b(N381), .out(\r126/LTV1 [57]) );
  nand2 \r126/ULTI1_57  ( .a(\r126/AEQB [57]), .b(\r126/LTV [57]), .out(
        \r126/LTV2 [57]) );
  nand2 \r126/ULTI2_57  ( .a(\r126/LTV1 [57]), .b(\r126/LTV2 [57]), .out(
        \r126/LTV [58]) );
  xor2 \r126/UEQI_58  ( .a(N444), .b(N380), .out(n2664) );
  nand2 \r126/UGTI0_58  ( .a(n2663), .b(N444), .out(\r126/GTV1 [58]) );
  nand2 \r126/UGTI1_58  ( .a(\r126/AEQB [58]), .b(\r126/GTV [58]), .out(
        \r126/GTV2 [58]) );
  nand2 \r126/UGTI2_58  ( .a(\r126/GTV1 [58]), .b(\r126/GTV2 [58]), .out(
        \r126/GTV [59]) );
  nand2 \r126/ULTI0_58  ( .a(n2662), .b(N380), .out(\r126/LTV1 [58]) );
  nand2 \r126/ULTI1_58  ( .a(\r126/AEQB [58]), .b(\r126/LTV [58]), .out(
        \r126/LTV2 [58]) );
  nand2 \r126/ULTI2_58  ( .a(\r126/LTV1 [58]), .b(\r126/LTV2 [58]), .out(
        \r126/LTV [59]) );
  xor2 \r126/UEQI_59  ( .a(N443), .b(N379), .out(n2661) );
  nand2 \r126/UGTI0_59  ( .a(n2660), .b(N443), .out(\r126/GTV1 [59]) );
  nand2 \r126/UGTI1_59  ( .a(\r126/AEQB [59]), .b(\r126/GTV [59]), .out(
        \r126/GTV2 [59]) );
  nand2 \r126/UGTI2_59  ( .a(\r126/GTV1 [59]), .b(\r126/GTV2 [59]), .out(
        \r126/GTV [60]) );
  nand2 \r126/ULTI0_59  ( .a(n2659), .b(N379), .out(\r126/LTV1 [59]) );
  nand2 \r126/ULTI1_59  ( .a(\r126/AEQB [59]), .b(\r126/LTV [59]), .out(
        \r126/LTV2 [59]) );
  nand2 \r126/ULTI2_59  ( .a(\r126/LTV1 [59]), .b(\r126/LTV2 [59]), .out(
        \r126/LTV [60]) );
  xor2 \r126/UEQI_60  ( .a(N442), .b(N378), .out(n2658) );
  nand2 \r126/UGTI0_60  ( .a(n2657), .b(N442), .out(\r126/GTV1 [60]) );
  nand2 \r126/UGTI1_60  ( .a(\r126/AEQB [60]), .b(\r126/GTV [60]), .out(
        \r126/GTV2 [60]) );
  nand2 \r126/UGTI2_60  ( .a(\r126/GTV1 [60]), .b(\r126/GTV2 [60]), .out(
        \r126/GTV [61]) );
  nand2 \r126/ULTI0_60  ( .a(n2656), .b(N378), .out(\r126/LTV1 [60]) );
  nand2 \r126/ULTI1_60  ( .a(\r126/AEQB [60]), .b(\r126/LTV [60]), .out(
        \r126/LTV2 [60]) );
  nand2 \r126/ULTI2_60  ( .a(\r126/LTV1 [60]), .b(\r126/LTV2 [60]), .out(
        \r126/LTV [61]) );
  xor2 \r126/UEQI_61  ( .a(N441), .b(N377), .out(n2655) );
  nand2 \r126/UGTI0_61  ( .a(n2654), .b(N441), .out(\r126/GTV1 [61]) );
  nand2 \r126/UGTI1_61  ( .a(\r126/AEQB [61]), .b(\r126/GTV [61]), .out(
        \r126/GTV2 [61]) );
  nand2 \r126/UGTI2_61  ( .a(\r126/GTV1 [61]), .b(\r126/GTV2 [61]), .out(
        \r126/GTV [62]) );
  nand2 \r126/ULTI0_61  ( .a(n2653), .b(N377), .out(\r126/LTV1 [61]) );
  nand2 \r126/ULTI1_61  ( .a(\r126/AEQB [61]), .b(\r126/LTV [61]), .out(
        \r126/LTV2 [61]) );
  nand2 \r126/ULTI2_61  ( .a(\r126/LTV1 [61]), .b(\r126/LTV2 [61]), .out(
        \r126/LTV [62]) );
  xor2 \r126/UEQI_62  ( .a(N440), .b(N376), .out(n2652) );
  nand2 \r126/UGTI0_62  ( .a(n2651), .b(N440), .out(\r126/GTV1 [62]) );
  nand2 \r126/UGTI1_62  ( .a(\r126/AEQB [62]), .b(\r126/GTV [62]), .out(
        \r126/GTV2 [62]) );
  nand2 \r126/UGTI2_62  ( .a(\r126/GTV1 [62]), .b(\r126/GTV2 [62]), .out(
        \r126/GTV [63]) );
  nand2 \r126/ULTI0_62  ( .a(n2650), .b(N376), .out(\r126/LTV1 [62]) );
  nand2 \r126/ULTI1_62  ( .a(\r126/AEQB [62]), .b(\r126/LTV [62]), .out(
        \r126/LTV2 [62]) );
  nand2 \r126/ULTI2_62  ( .a(\r126/LTV1 [62]), .b(\r126/LTV2 [62]), .out(
        \r126/LTV [63]) );
  nor2 \r125/UEQ  ( .a(N221), .b(N223), .out(N225) );
  nand2 \r125/UNGT0  ( .a(N218), .b(n2649), .out(n2648) );
  nand2 \r125/UNLT0  ( .a(N154), .b(n2647), .out(n2646) );
  xor2 \r125/UEQI  ( .a(\r125/SA ), .b(\r125/SB ), .out(n2645) );
  nand2 \r125/UGTI0  ( .a(n2644), .b(\r125/SA ), .out(\r125/GTV1 [63]) );
  nand2 \r125/UGTI1  ( .a(\r125/AEQB [63]), .b(\r125/GTV [63]), .out(
        \r125/GTV2 [63]) );
  nand2 \r125/UGTI2  ( .a(\r125/GTV1 [63]), .b(\r125/GTV2 [63]), .out(N221) );
  nand2 \r125/ULTI0  ( .a(n2643), .b(\r125/SB ), .out(\r125/LTV1 [63]) );
  nand2 \r125/ULTI1  ( .a(\r125/AEQB [63]), .b(\r125/LTV [63]), .out(
        \r125/LTV2 [63]) );
  nand2 \r125/ULTI2  ( .a(\r125/LTV1 [63]), .b(\r125/LTV2 [63]), .out(N223) );
  xor2 \r125/UEQI_1  ( .a(N217), .b(N153), .out(n2642) );
  nand2 \r125/UGTI0_1  ( .a(n2641), .b(N217), .out(\r125/GTV1 [1]) );
  nand2 \r125/UGTI1_1  ( .a(\r125/AEQB [1]), .b(\r125/GTV [1]), .out(
        \r125/GTV2 [1]) );
  nand2 \r125/UGTI2_1  ( .a(\r125/GTV1 [1]), .b(\r125/GTV2 [1]), .out(
        \r125/GTV [2]) );
  nand2 \r125/ULTI0_1  ( .a(n2640), .b(N153), .out(\r125/LTV1 [1]) );
  nand2 \r125/ULTI1_1  ( .a(\r125/AEQB [1]), .b(\r125/LTV [1]), .out(
        \r125/LTV2 [1]) );
  nand2 \r125/ULTI2_1  ( .a(\r125/LTV1 [1]), .b(\r125/LTV2 [1]), .out(
        \r125/LTV [2]) );
  xor2 \r125/UEQI_2  ( .a(N216), .b(N152), .out(n2639) );
  nand2 \r125/UGTI0_2  ( .a(n2638), .b(N216), .out(\r125/GTV1 [2]) );
  nand2 \r125/UGTI1_2  ( .a(\r125/AEQB [2]), .b(\r125/GTV [2]), .out(
        \r125/GTV2 [2]) );
  nand2 \r125/UGTI2_2  ( .a(\r125/GTV1 [2]), .b(\r125/GTV2 [2]), .out(
        \r125/GTV [3]) );
  nand2 \r125/ULTI0_2  ( .a(n2637), .b(N152), .out(\r125/LTV1 [2]) );
  nand2 \r125/ULTI1_2  ( .a(\r125/AEQB [2]), .b(\r125/LTV [2]), .out(
        \r125/LTV2 [2]) );
  nand2 \r125/ULTI2_2  ( .a(\r125/LTV1 [2]), .b(\r125/LTV2 [2]), .out(
        \r125/LTV [3]) );
  xor2 \r125/UEQI_3  ( .a(N215), .b(N151), .out(n2636) );
  nand2 \r125/UGTI0_3  ( .a(n2635), .b(N215), .out(\r125/GTV1 [3]) );
  nand2 \r125/UGTI1_3  ( .a(\r125/AEQB [3]), .b(\r125/GTV [3]), .out(
        \r125/GTV2 [3]) );
  nand2 \r125/UGTI2_3  ( .a(\r125/GTV1 [3]), .b(\r125/GTV2 [3]), .out(
        \r125/GTV [4]) );
  nand2 \r125/ULTI0_3  ( .a(n2634), .b(N151), .out(\r125/LTV1 [3]) );
  nand2 \r125/ULTI1_3  ( .a(\r125/AEQB [3]), .b(\r125/LTV [3]), .out(
        \r125/LTV2 [3]) );
  nand2 \r125/ULTI2_3  ( .a(\r125/LTV1 [3]), .b(\r125/LTV2 [3]), .out(
        \r125/LTV [4]) );
  xor2 \r125/UEQI_4  ( .a(N214), .b(N150), .out(n2633) );
  nand2 \r125/UGTI0_4  ( .a(n2632), .b(N214), .out(\r125/GTV1 [4]) );
  nand2 \r125/UGTI1_4  ( .a(\r125/AEQB [4]), .b(\r125/GTV [4]), .out(
        \r125/GTV2 [4]) );
  nand2 \r125/UGTI2_4  ( .a(\r125/GTV1 [4]), .b(\r125/GTV2 [4]), .out(
        \r125/GTV [5]) );
  nand2 \r125/ULTI0_4  ( .a(n2631), .b(N150), .out(\r125/LTV1 [4]) );
  nand2 \r125/ULTI1_4  ( .a(\r125/AEQB [4]), .b(\r125/LTV [4]), .out(
        \r125/LTV2 [4]) );
  nand2 \r125/ULTI2_4  ( .a(\r125/LTV1 [4]), .b(\r125/LTV2 [4]), .out(
        \r125/LTV [5]) );
  xor2 \r125/UEQI_5  ( .a(N213), .b(N149), .out(n2630) );
  nand2 \r125/UGTI0_5  ( .a(n2629), .b(N213), .out(\r125/GTV1 [5]) );
  nand2 \r125/UGTI1_5  ( .a(\r125/AEQB [5]), .b(\r125/GTV [5]), .out(
        \r125/GTV2 [5]) );
  nand2 \r125/UGTI2_5  ( .a(\r125/GTV1 [5]), .b(\r125/GTV2 [5]), .out(
        \r125/GTV [6]) );
  nand2 \r125/ULTI0_5  ( .a(n2628), .b(N149), .out(\r125/LTV1 [5]) );
  nand2 \r125/ULTI1_5  ( .a(\r125/AEQB [5]), .b(\r125/LTV [5]), .out(
        \r125/LTV2 [5]) );
  nand2 \r125/ULTI2_5  ( .a(\r125/LTV1 [5]), .b(\r125/LTV2 [5]), .out(
        \r125/LTV [6]) );
  xor2 \r125/UEQI_6  ( .a(N212), .b(N148), .out(n2627) );
  nand2 \r125/UGTI0_6  ( .a(n2626), .b(N212), .out(\r125/GTV1 [6]) );
  nand2 \r125/UGTI1_6  ( .a(\r125/AEQB [6]), .b(\r125/GTV [6]), .out(
        \r125/GTV2 [6]) );
  nand2 \r125/UGTI2_6  ( .a(\r125/GTV1 [6]), .b(\r125/GTV2 [6]), .out(
        \r125/GTV [7]) );
  nand2 \r125/ULTI0_6  ( .a(n2625), .b(N148), .out(\r125/LTV1 [6]) );
  nand2 \r125/ULTI1_6  ( .a(\r125/AEQB [6]), .b(\r125/LTV [6]), .out(
        \r125/LTV2 [6]) );
  nand2 \r125/ULTI2_6  ( .a(\r125/LTV1 [6]), .b(\r125/LTV2 [6]), .out(
        \r125/LTV [7]) );
  xor2 \r125/UEQI_7  ( .a(N211), .b(N147), .out(n2624) );
  nand2 \r125/UGTI0_7  ( .a(n2623), .b(N211), .out(\r125/GTV1 [7]) );
  nand2 \r125/UGTI1_7  ( .a(\r125/AEQB [7]), .b(\r125/GTV [7]), .out(
        \r125/GTV2 [7]) );
  nand2 \r125/UGTI2_7  ( .a(\r125/GTV1 [7]), .b(\r125/GTV2 [7]), .out(
        \r125/GTV [8]) );
  nand2 \r125/ULTI0_7  ( .a(n2622), .b(N147), .out(\r125/LTV1 [7]) );
  nand2 \r125/ULTI1_7  ( .a(\r125/AEQB [7]), .b(\r125/LTV [7]), .out(
        \r125/LTV2 [7]) );
  nand2 \r125/ULTI2_7  ( .a(\r125/LTV1 [7]), .b(\r125/LTV2 [7]), .out(
        \r125/LTV [8]) );
  xor2 \r125/UEQI_8  ( .a(N210), .b(N146), .out(n2621) );
  nand2 \r125/UGTI0_8  ( .a(n2620), .b(N210), .out(\r125/GTV1 [8]) );
  nand2 \r125/UGTI1_8  ( .a(\r125/AEQB [8]), .b(\r125/GTV [8]), .out(
        \r125/GTV2 [8]) );
  nand2 \r125/UGTI2_8  ( .a(\r125/GTV1 [8]), .b(\r125/GTV2 [8]), .out(
        \r125/GTV [9]) );
  nand2 \r125/ULTI0_8  ( .a(n2619), .b(N146), .out(\r125/LTV1 [8]) );
  nand2 \r125/ULTI1_8  ( .a(\r125/AEQB [8]), .b(\r125/LTV [8]), .out(
        \r125/LTV2 [8]) );
  nand2 \r125/ULTI2_8  ( .a(\r125/LTV1 [8]), .b(\r125/LTV2 [8]), .out(
        \r125/LTV [9]) );
  xor2 \r125/UEQI_9  ( .a(N209), .b(N145), .out(n2618) );
  nand2 \r125/UGTI0_9  ( .a(n2617), .b(N209), .out(\r125/GTV1 [9]) );
  nand2 \r125/UGTI1_9  ( .a(\r125/AEQB [9]), .b(\r125/GTV [9]), .out(
        \r125/GTV2 [9]) );
  nand2 \r125/UGTI2_9  ( .a(\r125/GTV1 [9]), .b(\r125/GTV2 [9]), .out(
        \r125/GTV [10]) );
  nand2 \r125/ULTI0_9  ( .a(n2616), .b(N145), .out(\r125/LTV1 [9]) );
  nand2 \r125/ULTI1_9  ( .a(\r125/AEQB [9]), .b(\r125/LTV [9]), .out(
        \r125/LTV2 [9]) );
  nand2 \r125/ULTI2_9  ( .a(\r125/LTV1 [9]), .b(\r125/LTV2 [9]), .out(
        \r125/LTV [10]) );
  xor2 \r125/UEQI_10  ( .a(N208), .b(N144), .out(n2615) );
  nand2 \r125/UGTI0_10  ( .a(n2614), .b(N208), .out(\r125/GTV1 [10]) );
  nand2 \r125/UGTI1_10  ( .a(\r125/AEQB [10]), .b(\r125/GTV [10]), .out(
        \r125/GTV2 [10]) );
  nand2 \r125/UGTI2_10  ( .a(\r125/GTV1 [10]), .b(\r125/GTV2 [10]), .out(
        \r125/GTV [11]) );
  nand2 \r125/ULTI0_10  ( .a(n2613), .b(N144), .out(\r125/LTV1 [10]) );
  nand2 \r125/ULTI1_10  ( .a(\r125/AEQB [10]), .b(\r125/LTV [10]), .out(
        \r125/LTV2 [10]) );
  nand2 \r125/ULTI2_10  ( .a(\r125/LTV1 [10]), .b(\r125/LTV2 [10]), .out(
        \r125/LTV [11]) );
  xor2 \r125/UEQI_11  ( .a(N207), .b(N143), .out(n2612) );
  nand2 \r125/UGTI0_11  ( .a(n2611), .b(N207), .out(\r125/GTV1 [11]) );
  nand2 \r125/UGTI1_11  ( .a(\r125/AEQB [11]), .b(\r125/GTV [11]), .out(
        \r125/GTV2 [11]) );
  nand2 \r125/UGTI2_11  ( .a(\r125/GTV1 [11]), .b(\r125/GTV2 [11]), .out(
        \r125/GTV [12]) );
  nand2 \r125/ULTI0_11  ( .a(n2610), .b(N143), .out(\r125/LTV1 [11]) );
  nand2 \r125/ULTI1_11  ( .a(\r125/AEQB [11]), .b(\r125/LTV [11]), .out(
        \r125/LTV2 [11]) );
  nand2 \r125/ULTI2_11  ( .a(\r125/LTV1 [11]), .b(\r125/LTV2 [11]), .out(
        \r125/LTV [12]) );
  xor2 \r125/UEQI_12  ( .a(N206), .b(N142), .out(n2609) );
  nand2 \r125/UGTI0_12  ( .a(n2608), .b(N206), .out(\r125/GTV1 [12]) );
  nand2 \r125/UGTI1_12  ( .a(\r125/AEQB [12]), .b(\r125/GTV [12]), .out(
        \r125/GTV2 [12]) );
  nand2 \r125/UGTI2_12  ( .a(\r125/GTV1 [12]), .b(\r125/GTV2 [12]), .out(
        \r125/GTV [13]) );
  nand2 \r125/ULTI0_12  ( .a(n2607), .b(N142), .out(\r125/LTV1 [12]) );
  nand2 \r125/ULTI1_12  ( .a(\r125/AEQB [12]), .b(\r125/LTV [12]), .out(
        \r125/LTV2 [12]) );
  nand2 \r125/ULTI2_12  ( .a(\r125/LTV1 [12]), .b(\r125/LTV2 [12]), .out(
        \r125/LTV [13]) );
  xor2 \r125/UEQI_13  ( .a(N205), .b(N141), .out(n2606) );
  nand2 \r125/UGTI0_13  ( .a(n2605), .b(N205), .out(\r125/GTV1 [13]) );
  nand2 \r125/UGTI1_13  ( .a(\r125/AEQB [13]), .b(\r125/GTV [13]), .out(
        \r125/GTV2 [13]) );
  nand2 \r125/UGTI2_13  ( .a(\r125/GTV1 [13]), .b(\r125/GTV2 [13]), .out(
        \r125/GTV [14]) );
  nand2 \r125/ULTI0_13  ( .a(n2604), .b(N141), .out(\r125/LTV1 [13]) );
  nand2 \r125/ULTI1_13  ( .a(\r125/AEQB [13]), .b(\r125/LTV [13]), .out(
        \r125/LTV2 [13]) );
  nand2 \r125/ULTI2_13  ( .a(\r125/LTV1 [13]), .b(\r125/LTV2 [13]), .out(
        \r125/LTV [14]) );
  xor2 \r125/UEQI_14  ( .a(N204), .b(N140), .out(n2603) );
  nand2 \r125/UGTI0_14  ( .a(n2602), .b(N204), .out(\r125/GTV1 [14]) );
  nand2 \r125/UGTI1_14  ( .a(\r125/AEQB [14]), .b(\r125/GTV [14]), .out(
        \r125/GTV2 [14]) );
  nand2 \r125/UGTI2_14  ( .a(\r125/GTV1 [14]), .b(\r125/GTV2 [14]), .out(
        \r125/GTV [15]) );
  nand2 \r125/ULTI0_14  ( .a(n2601), .b(N140), .out(\r125/LTV1 [14]) );
  nand2 \r125/ULTI1_14  ( .a(\r125/AEQB [14]), .b(\r125/LTV [14]), .out(
        \r125/LTV2 [14]) );
  nand2 \r125/ULTI2_14  ( .a(\r125/LTV1 [14]), .b(\r125/LTV2 [14]), .out(
        \r125/LTV [15]) );
  xor2 \r125/UEQI_15  ( .a(N203), .b(N139), .out(n2600) );
  nand2 \r125/UGTI0_15  ( .a(n2599), .b(N203), .out(\r125/GTV1 [15]) );
  nand2 \r125/UGTI1_15  ( .a(\r125/AEQB [15]), .b(\r125/GTV [15]), .out(
        \r125/GTV2 [15]) );
  nand2 \r125/UGTI2_15  ( .a(\r125/GTV1 [15]), .b(\r125/GTV2 [15]), .out(
        \r125/GTV [16]) );
  nand2 \r125/ULTI0_15  ( .a(n2598), .b(N139), .out(\r125/LTV1 [15]) );
  nand2 \r125/ULTI1_15  ( .a(\r125/AEQB [15]), .b(\r125/LTV [15]), .out(
        \r125/LTV2 [15]) );
  nand2 \r125/ULTI2_15  ( .a(\r125/LTV1 [15]), .b(\r125/LTV2 [15]), .out(
        \r125/LTV [16]) );
  xor2 \r125/UEQI_16  ( .a(N202), .b(N138), .out(n2597) );
  nand2 \r125/UGTI0_16  ( .a(n2596), .b(N202), .out(\r125/GTV1 [16]) );
  nand2 \r125/UGTI1_16  ( .a(\r125/AEQB [16]), .b(\r125/GTV [16]), .out(
        \r125/GTV2 [16]) );
  nand2 \r125/UGTI2_16  ( .a(\r125/GTV1 [16]), .b(\r125/GTV2 [16]), .out(
        \r125/GTV [17]) );
  nand2 \r125/ULTI0_16  ( .a(n2595), .b(N138), .out(\r125/LTV1 [16]) );
  nand2 \r125/ULTI1_16  ( .a(\r125/AEQB [16]), .b(\r125/LTV [16]), .out(
        \r125/LTV2 [16]) );
  nand2 \r125/ULTI2_16  ( .a(\r125/LTV1 [16]), .b(\r125/LTV2 [16]), .out(
        \r125/LTV [17]) );
  xor2 \r125/UEQI_17  ( .a(N201), .b(N137), .out(n2594) );
  nand2 \r125/UGTI0_17  ( .a(n2593), .b(N201), .out(\r125/GTV1 [17]) );
  nand2 \r125/UGTI1_17  ( .a(\r125/AEQB [17]), .b(\r125/GTV [17]), .out(
        \r125/GTV2 [17]) );
  nand2 \r125/UGTI2_17  ( .a(\r125/GTV1 [17]), .b(\r125/GTV2 [17]), .out(
        \r125/GTV [18]) );
  nand2 \r125/ULTI0_17  ( .a(n2592), .b(N137), .out(\r125/LTV1 [17]) );
  nand2 \r125/ULTI1_17  ( .a(\r125/AEQB [17]), .b(\r125/LTV [17]), .out(
        \r125/LTV2 [17]) );
  nand2 \r125/ULTI2_17  ( .a(\r125/LTV1 [17]), .b(\r125/LTV2 [17]), .out(
        \r125/LTV [18]) );
  xor2 \r125/UEQI_18  ( .a(N200), .b(N136), .out(n2591) );
  nand2 \r125/UGTI0_18  ( .a(n2590), .b(N200), .out(\r125/GTV1 [18]) );
  nand2 \r125/UGTI1_18  ( .a(\r125/AEQB [18]), .b(\r125/GTV [18]), .out(
        \r125/GTV2 [18]) );
  nand2 \r125/UGTI2_18  ( .a(\r125/GTV1 [18]), .b(\r125/GTV2 [18]), .out(
        \r125/GTV [19]) );
  nand2 \r125/ULTI0_18  ( .a(n2589), .b(N136), .out(\r125/LTV1 [18]) );
  nand2 \r125/ULTI1_18  ( .a(\r125/AEQB [18]), .b(\r125/LTV [18]), .out(
        \r125/LTV2 [18]) );
  nand2 \r125/ULTI2_18  ( .a(\r125/LTV1 [18]), .b(\r125/LTV2 [18]), .out(
        \r125/LTV [19]) );
  xor2 \r125/UEQI_19  ( .a(N199), .b(N135), .out(n2588) );
  nand2 \r125/UGTI0_19  ( .a(n2587), .b(N199), .out(\r125/GTV1 [19]) );
  nand2 \r125/UGTI1_19  ( .a(\r125/AEQB [19]), .b(\r125/GTV [19]), .out(
        \r125/GTV2 [19]) );
  nand2 \r125/UGTI2_19  ( .a(\r125/GTV1 [19]), .b(\r125/GTV2 [19]), .out(
        \r125/GTV [20]) );
  nand2 \r125/ULTI0_19  ( .a(n2586), .b(N135), .out(\r125/LTV1 [19]) );
  nand2 \r125/ULTI1_19  ( .a(\r125/AEQB [19]), .b(\r125/LTV [19]), .out(
        \r125/LTV2 [19]) );
  nand2 \r125/ULTI2_19  ( .a(\r125/LTV1 [19]), .b(\r125/LTV2 [19]), .out(
        \r125/LTV [20]) );
  xor2 \r125/UEQI_20  ( .a(N198), .b(N134), .out(n2585) );
  nand2 \r125/UGTI0_20  ( .a(n2584), .b(N198), .out(\r125/GTV1 [20]) );
  nand2 \r125/UGTI1_20  ( .a(\r125/AEQB [20]), .b(\r125/GTV [20]), .out(
        \r125/GTV2 [20]) );
  nand2 \r125/UGTI2_20  ( .a(\r125/GTV1 [20]), .b(\r125/GTV2 [20]), .out(
        \r125/GTV [21]) );
  nand2 \r125/ULTI0_20  ( .a(n2583), .b(N134), .out(\r125/LTV1 [20]) );
  nand2 \r125/ULTI1_20  ( .a(\r125/AEQB [20]), .b(\r125/LTV [20]), .out(
        \r125/LTV2 [20]) );
  nand2 \r125/ULTI2_20  ( .a(\r125/LTV1 [20]), .b(\r125/LTV2 [20]), .out(
        \r125/LTV [21]) );
  xor2 \r125/UEQI_21  ( .a(N197), .b(N133), .out(n2582) );
  nand2 \r125/UGTI0_21  ( .a(n2581), .b(N197), .out(\r125/GTV1 [21]) );
  nand2 \r125/UGTI1_21  ( .a(\r125/AEQB [21]), .b(\r125/GTV [21]), .out(
        \r125/GTV2 [21]) );
  nand2 \r125/UGTI2_21  ( .a(\r125/GTV1 [21]), .b(\r125/GTV2 [21]), .out(
        \r125/GTV [22]) );
  nand2 \r125/ULTI0_21  ( .a(n2580), .b(N133), .out(\r125/LTV1 [21]) );
  nand2 \r125/ULTI1_21  ( .a(\r125/AEQB [21]), .b(\r125/LTV [21]), .out(
        \r125/LTV2 [21]) );
  nand2 \r125/ULTI2_21  ( .a(\r125/LTV1 [21]), .b(\r125/LTV2 [21]), .out(
        \r125/LTV [22]) );
  xor2 \r125/UEQI_22  ( .a(N196), .b(N132), .out(n2579) );
  nand2 \r125/UGTI0_22  ( .a(n2578), .b(N196), .out(\r125/GTV1 [22]) );
  nand2 \r125/UGTI1_22  ( .a(\r125/AEQB [22]), .b(\r125/GTV [22]), .out(
        \r125/GTV2 [22]) );
  nand2 \r125/UGTI2_22  ( .a(\r125/GTV1 [22]), .b(\r125/GTV2 [22]), .out(
        \r125/GTV [23]) );
  nand2 \r125/ULTI0_22  ( .a(n2577), .b(N132), .out(\r125/LTV1 [22]) );
  nand2 \r125/ULTI1_22  ( .a(\r125/AEQB [22]), .b(\r125/LTV [22]), .out(
        \r125/LTV2 [22]) );
  nand2 \r125/ULTI2_22  ( .a(\r125/LTV1 [22]), .b(\r125/LTV2 [22]), .out(
        \r125/LTV [23]) );
  xor2 \r125/UEQI_23  ( .a(N195), .b(N131), .out(n2576) );
  nand2 \r125/UGTI0_23  ( .a(n2575), .b(N195), .out(\r125/GTV1 [23]) );
  nand2 \r125/UGTI1_23  ( .a(\r125/AEQB [23]), .b(\r125/GTV [23]), .out(
        \r125/GTV2 [23]) );
  nand2 \r125/UGTI2_23  ( .a(\r125/GTV1 [23]), .b(\r125/GTV2 [23]), .out(
        \r125/GTV [24]) );
  nand2 \r125/ULTI0_23  ( .a(n2574), .b(N131), .out(\r125/LTV1 [23]) );
  nand2 \r125/ULTI1_23  ( .a(\r125/AEQB [23]), .b(\r125/LTV [23]), .out(
        \r125/LTV2 [23]) );
  nand2 \r125/ULTI2_23  ( .a(\r125/LTV1 [23]), .b(\r125/LTV2 [23]), .out(
        \r125/LTV [24]) );
  xor2 \r125/UEQI_24  ( .a(N194), .b(N130), .out(n2573) );
  nand2 \r125/UGTI0_24  ( .a(n2572), .b(N194), .out(\r125/GTV1 [24]) );
  nand2 \r125/UGTI1_24  ( .a(\r125/AEQB [24]), .b(\r125/GTV [24]), .out(
        \r125/GTV2 [24]) );
  nand2 \r125/UGTI2_24  ( .a(\r125/GTV1 [24]), .b(\r125/GTV2 [24]), .out(
        \r125/GTV [25]) );
  nand2 \r125/ULTI0_24  ( .a(n2571), .b(N130), .out(\r125/LTV1 [24]) );
  nand2 \r125/ULTI1_24  ( .a(\r125/AEQB [24]), .b(\r125/LTV [24]), .out(
        \r125/LTV2 [24]) );
  nand2 \r125/ULTI2_24  ( .a(\r125/LTV1 [24]), .b(\r125/LTV2 [24]), .out(
        \r125/LTV [25]) );
  xor2 \r125/UEQI_25  ( .a(N193), .b(N129), .out(n2570) );
  nand2 \r125/UGTI0_25  ( .a(n2569), .b(N193), .out(\r125/GTV1 [25]) );
  nand2 \r125/UGTI1_25  ( .a(\r125/AEQB [25]), .b(\r125/GTV [25]), .out(
        \r125/GTV2 [25]) );
  nand2 \r125/UGTI2_25  ( .a(\r125/GTV1 [25]), .b(\r125/GTV2 [25]), .out(
        \r125/GTV [26]) );
  nand2 \r125/ULTI0_25  ( .a(n2568), .b(N129), .out(\r125/LTV1 [25]) );
  nand2 \r125/ULTI1_25  ( .a(\r125/AEQB [25]), .b(\r125/LTV [25]), .out(
        \r125/LTV2 [25]) );
  nand2 \r125/ULTI2_25  ( .a(\r125/LTV1 [25]), .b(\r125/LTV2 [25]), .out(
        \r125/LTV [26]) );
  xor2 \r125/UEQI_26  ( .a(N192), .b(N128), .out(n2567) );
  nand2 \r125/UGTI0_26  ( .a(n2566), .b(N192), .out(\r125/GTV1 [26]) );
  nand2 \r125/UGTI1_26  ( .a(\r125/AEQB [26]), .b(\r125/GTV [26]), .out(
        \r125/GTV2 [26]) );
  nand2 \r125/UGTI2_26  ( .a(\r125/GTV1 [26]), .b(\r125/GTV2 [26]), .out(
        \r125/GTV [27]) );
  nand2 \r125/ULTI0_26  ( .a(n2565), .b(N128), .out(\r125/LTV1 [26]) );
  nand2 \r125/ULTI1_26  ( .a(\r125/AEQB [26]), .b(\r125/LTV [26]), .out(
        \r125/LTV2 [26]) );
  nand2 \r125/ULTI2_26  ( .a(\r125/LTV1 [26]), .b(\r125/LTV2 [26]), .out(
        \r125/LTV [27]) );
  xor2 \r125/UEQI_27  ( .a(N191), .b(N127), .out(n2564) );
  nand2 \r125/UGTI0_27  ( .a(n2563), .b(N191), .out(\r125/GTV1 [27]) );
  nand2 \r125/UGTI1_27  ( .a(\r125/AEQB [27]), .b(\r125/GTV [27]), .out(
        \r125/GTV2 [27]) );
  nand2 \r125/UGTI2_27  ( .a(\r125/GTV1 [27]), .b(\r125/GTV2 [27]), .out(
        \r125/GTV [28]) );
  nand2 \r125/ULTI0_27  ( .a(n2562), .b(N127), .out(\r125/LTV1 [27]) );
  nand2 \r125/ULTI1_27  ( .a(\r125/AEQB [27]), .b(\r125/LTV [27]), .out(
        \r125/LTV2 [27]) );
  nand2 \r125/ULTI2_27  ( .a(\r125/LTV1 [27]), .b(\r125/LTV2 [27]), .out(
        \r125/LTV [28]) );
  xor2 \r125/UEQI_28  ( .a(N190), .b(N126), .out(n2561) );
  nand2 \r125/UGTI0_28  ( .a(n2560), .b(N190), .out(\r125/GTV1 [28]) );
  nand2 \r125/UGTI1_28  ( .a(\r125/AEQB [28]), .b(\r125/GTV [28]), .out(
        \r125/GTV2 [28]) );
  nand2 \r125/UGTI2_28  ( .a(\r125/GTV1 [28]), .b(\r125/GTV2 [28]), .out(
        \r125/GTV [29]) );
  nand2 \r125/ULTI0_28  ( .a(n2559), .b(N126), .out(\r125/LTV1 [28]) );
  nand2 \r125/ULTI1_28  ( .a(\r125/AEQB [28]), .b(\r125/LTV [28]), .out(
        \r125/LTV2 [28]) );
  nand2 \r125/ULTI2_28  ( .a(\r125/LTV1 [28]), .b(\r125/LTV2 [28]), .out(
        \r125/LTV [29]) );
  xor2 \r125/UEQI_29  ( .a(N189), .b(N125), .out(n2558) );
  nand2 \r125/UGTI0_29  ( .a(n2557), .b(N189), .out(\r125/GTV1 [29]) );
  nand2 \r125/UGTI1_29  ( .a(\r125/AEQB [29]), .b(\r125/GTV [29]), .out(
        \r125/GTV2 [29]) );
  nand2 \r125/UGTI2_29  ( .a(\r125/GTV1 [29]), .b(\r125/GTV2 [29]), .out(
        \r125/GTV [30]) );
  nand2 \r125/ULTI0_29  ( .a(n2556), .b(N125), .out(\r125/LTV1 [29]) );
  nand2 \r125/ULTI1_29  ( .a(\r125/AEQB [29]), .b(\r125/LTV [29]), .out(
        \r125/LTV2 [29]) );
  nand2 \r125/ULTI2_29  ( .a(\r125/LTV1 [29]), .b(\r125/LTV2 [29]), .out(
        \r125/LTV [30]) );
  xor2 \r125/UEQI_30  ( .a(N188), .b(N124), .out(n2555) );
  nand2 \r125/UGTI0_30  ( .a(n2554), .b(N188), .out(\r125/GTV1 [30]) );
  nand2 \r125/UGTI1_30  ( .a(\r125/AEQB [30]), .b(\r125/GTV [30]), .out(
        \r125/GTV2 [30]) );
  nand2 \r125/UGTI2_30  ( .a(\r125/GTV1 [30]), .b(\r125/GTV2 [30]), .out(
        \r125/GTV [31]) );
  nand2 \r125/ULTI0_30  ( .a(n2553), .b(N124), .out(\r125/LTV1 [30]) );
  nand2 \r125/ULTI1_30  ( .a(\r125/AEQB [30]), .b(\r125/LTV [30]), .out(
        \r125/LTV2 [30]) );
  nand2 \r125/ULTI2_30  ( .a(\r125/LTV1 [30]), .b(\r125/LTV2 [30]), .out(
        \r125/LTV [31]) );
  xor2 \r125/UEQI_31  ( .a(N187), .b(N123), .out(n2552) );
  nand2 \r125/UGTI0_31  ( .a(n2551), .b(N187), .out(\r125/GTV1 [31]) );
  nand2 \r125/UGTI1_31  ( .a(\r125/AEQB [31]), .b(\r125/GTV [31]), .out(
        \r125/GTV2 [31]) );
  nand2 \r125/UGTI2_31  ( .a(\r125/GTV1 [31]), .b(\r125/GTV2 [31]), .out(
        \r125/GTV [32]) );
  nand2 \r125/ULTI0_31  ( .a(n2550), .b(N123), .out(\r125/LTV1 [31]) );
  nand2 \r125/ULTI1_31  ( .a(\r125/AEQB [31]), .b(\r125/LTV [31]), .out(
        \r125/LTV2 [31]) );
  nand2 \r125/ULTI2_31  ( .a(\r125/LTV1 [31]), .b(\r125/LTV2 [31]), .out(
        \r125/LTV [32]) );
  xor2 \r125/UEQI_32  ( .a(N186), .b(N122), .out(n2549) );
  nand2 \r125/UGTI0_32  ( .a(n2548), .b(N186), .out(\r125/GTV1 [32]) );
  nand2 \r125/UGTI1_32  ( .a(\r125/AEQB [32]), .b(\r125/GTV [32]), .out(
        \r125/GTV2 [32]) );
  nand2 \r125/UGTI2_32  ( .a(\r125/GTV1 [32]), .b(\r125/GTV2 [32]), .out(
        \r125/GTV [33]) );
  nand2 \r125/ULTI0_32  ( .a(n2547), .b(N122), .out(\r125/LTV1 [32]) );
  nand2 \r125/ULTI1_32  ( .a(\r125/AEQB [32]), .b(\r125/LTV [32]), .out(
        \r125/LTV2 [32]) );
  nand2 \r125/ULTI2_32  ( .a(\r125/LTV1 [32]), .b(\r125/LTV2 [32]), .out(
        \r125/LTV [33]) );
  xor2 \r125/UEQI_33  ( .a(N185), .b(N121), .out(n2546) );
  nand2 \r125/UGTI0_33  ( .a(n2545), .b(N185), .out(\r125/GTV1 [33]) );
  nand2 \r125/UGTI1_33  ( .a(\r125/AEQB [33]), .b(\r125/GTV [33]), .out(
        \r125/GTV2 [33]) );
  nand2 \r125/UGTI2_33  ( .a(\r125/GTV1 [33]), .b(\r125/GTV2 [33]), .out(
        \r125/GTV [34]) );
  nand2 \r125/ULTI0_33  ( .a(n2544), .b(N121), .out(\r125/LTV1 [33]) );
  nand2 \r125/ULTI1_33  ( .a(\r125/AEQB [33]), .b(\r125/LTV [33]), .out(
        \r125/LTV2 [33]) );
  nand2 \r125/ULTI2_33  ( .a(\r125/LTV1 [33]), .b(\r125/LTV2 [33]), .out(
        \r125/LTV [34]) );
  xor2 \r125/UEQI_34  ( .a(N184), .b(N120), .out(n2543) );
  nand2 \r125/UGTI0_34  ( .a(n2542), .b(N184), .out(\r125/GTV1 [34]) );
  nand2 \r125/UGTI1_34  ( .a(\r125/AEQB [34]), .b(\r125/GTV [34]), .out(
        \r125/GTV2 [34]) );
  nand2 \r125/UGTI2_34  ( .a(\r125/GTV1 [34]), .b(\r125/GTV2 [34]), .out(
        \r125/GTV [35]) );
  nand2 \r125/ULTI0_34  ( .a(n2541), .b(N120), .out(\r125/LTV1 [34]) );
  nand2 \r125/ULTI1_34  ( .a(\r125/AEQB [34]), .b(\r125/LTV [34]), .out(
        \r125/LTV2 [34]) );
  nand2 \r125/ULTI2_34  ( .a(\r125/LTV1 [34]), .b(\r125/LTV2 [34]), .out(
        \r125/LTV [35]) );
  xor2 \r125/UEQI_35  ( .a(N183), .b(N119), .out(n2540) );
  nand2 \r125/UGTI0_35  ( .a(n2539), .b(N183), .out(\r125/GTV1 [35]) );
  nand2 \r125/UGTI1_35  ( .a(\r125/AEQB [35]), .b(\r125/GTV [35]), .out(
        \r125/GTV2 [35]) );
  nand2 \r125/UGTI2_35  ( .a(\r125/GTV1 [35]), .b(\r125/GTV2 [35]), .out(
        \r125/GTV [36]) );
  nand2 \r125/ULTI0_35  ( .a(n2538), .b(N119), .out(\r125/LTV1 [35]) );
  nand2 \r125/ULTI1_35  ( .a(\r125/AEQB [35]), .b(\r125/LTV [35]), .out(
        \r125/LTV2 [35]) );
  nand2 \r125/ULTI2_35  ( .a(\r125/LTV1 [35]), .b(\r125/LTV2 [35]), .out(
        \r125/LTV [36]) );
  xor2 \r125/UEQI_36  ( .a(N182), .b(N118), .out(n2537) );
  nand2 \r125/UGTI0_36  ( .a(n2536), .b(N182), .out(\r125/GTV1 [36]) );
  nand2 \r125/UGTI1_36  ( .a(\r125/AEQB [36]), .b(\r125/GTV [36]), .out(
        \r125/GTV2 [36]) );
  nand2 \r125/UGTI2_36  ( .a(\r125/GTV1 [36]), .b(\r125/GTV2 [36]), .out(
        \r125/GTV [37]) );
  nand2 \r125/ULTI0_36  ( .a(n2535), .b(N118), .out(\r125/LTV1 [36]) );
  nand2 \r125/ULTI1_36  ( .a(\r125/AEQB [36]), .b(\r125/LTV [36]), .out(
        \r125/LTV2 [36]) );
  nand2 \r125/ULTI2_36  ( .a(\r125/LTV1 [36]), .b(\r125/LTV2 [36]), .out(
        \r125/LTV [37]) );
  xor2 \r125/UEQI_37  ( .a(N181), .b(N117), .out(n2534) );
  nand2 \r125/UGTI0_37  ( .a(n2533), .b(N181), .out(\r125/GTV1 [37]) );
  nand2 \r125/UGTI1_37  ( .a(\r125/AEQB [37]), .b(\r125/GTV [37]), .out(
        \r125/GTV2 [37]) );
  nand2 \r125/UGTI2_37  ( .a(\r125/GTV1 [37]), .b(\r125/GTV2 [37]), .out(
        \r125/GTV [38]) );
  nand2 \r125/ULTI0_37  ( .a(n2532), .b(N117), .out(\r125/LTV1 [37]) );
  nand2 \r125/ULTI1_37  ( .a(\r125/AEQB [37]), .b(\r125/LTV [37]), .out(
        \r125/LTV2 [37]) );
  nand2 \r125/ULTI2_37  ( .a(\r125/LTV1 [37]), .b(\r125/LTV2 [37]), .out(
        \r125/LTV [38]) );
  xor2 \r125/UEQI_38  ( .a(N180), .b(N116), .out(n2531) );
  nand2 \r125/UGTI0_38  ( .a(n2530), .b(N180), .out(\r125/GTV1 [38]) );
  nand2 \r125/UGTI1_38  ( .a(\r125/AEQB [38]), .b(\r125/GTV [38]), .out(
        \r125/GTV2 [38]) );
  nand2 \r125/UGTI2_38  ( .a(\r125/GTV1 [38]), .b(\r125/GTV2 [38]), .out(
        \r125/GTV [39]) );
  nand2 \r125/ULTI0_38  ( .a(n2529), .b(N116), .out(\r125/LTV1 [38]) );
  nand2 \r125/ULTI1_38  ( .a(\r125/AEQB [38]), .b(\r125/LTV [38]), .out(
        \r125/LTV2 [38]) );
  nand2 \r125/ULTI2_38  ( .a(\r125/LTV1 [38]), .b(\r125/LTV2 [38]), .out(
        \r125/LTV [39]) );
  xor2 \r125/UEQI_39  ( .a(N179), .b(N115), .out(n2528) );
  nand2 \r125/UGTI0_39  ( .a(n2527), .b(N179), .out(\r125/GTV1 [39]) );
  nand2 \r125/UGTI1_39  ( .a(\r125/AEQB [39]), .b(\r125/GTV [39]), .out(
        \r125/GTV2 [39]) );
  nand2 \r125/UGTI2_39  ( .a(\r125/GTV1 [39]), .b(\r125/GTV2 [39]), .out(
        \r125/GTV [40]) );
  nand2 \r125/ULTI0_39  ( .a(n2526), .b(N115), .out(\r125/LTV1 [39]) );
  nand2 \r125/ULTI1_39  ( .a(\r125/AEQB [39]), .b(\r125/LTV [39]), .out(
        \r125/LTV2 [39]) );
  nand2 \r125/ULTI2_39  ( .a(\r125/LTV1 [39]), .b(\r125/LTV2 [39]), .out(
        \r125/LTV [40]) );
  xor2 \r125/UEQI_40  ( .a(N178), .b(N114), .out(n2525) );
  nand2 \r125/UGTI0_40  ( .a(n2524), .b(N178), .out(\r125/GTV1 [40]) );
  nand2 \r125/UGTI1_40  ( .a(\r125/AEQB [40]), .b(\r125/GTV [40]), .out(
        \r125/GTV2 [40]) );
  nand2 \r125/UGTI2_40  ( .a(\r125/GTV1 [40]), .b(\r125/GTV2 [40]), .out(
        \r125/GTV [41]) );
  nand2 \r125/ULTI0_40  ( .a(n2523), .b(N114), .out(\r125/LTV1 [40]) );
  nand2 \r125/ULTI1_40  ( .a(\r125/AEQB [40]), .b(\r125/LTV [40]), .out(
        \r125/LTV2 [40]) );
  nand2 \r125/ULTI2_40  ( .a(\r125/LTV1 [40]), .b(\r125/LTV2 [40]), .out(
        \r125/LTV [41]) );
  xor2 \r125/UEQI_41  ( .a(N177), .b(N113), .out(n2522) );
  nand2 \r125/UGTI0_41  ( .a(n2521), .b(N177), .out(\r125/GTV1 [41]) );
  nand2 \r125/UGTI1_41  ( .a(\r125/AEQB [41]), .b(\r125/GTV [41]), .out(
        \r125/GTV2 [41]) );
  nand2 \r125/UGTI2_41  ( .a(\r125/GTV1 [41]), .b(\r125/GTV2 [41]), .out(
        \r125/GTV [42]) );
  nand2 \r125/ULTI0_41  ( .a(n2520), .b(N113), .out(\r125/LTV1 [41]) );
  nand2 \r125/ULTI1_41  ( .a(\r125/AEQB [41]), .b(\r125/LTV [41]), .out(
        \r125/LTV2 [41]) );
  nand2 \r125/ULTI2_41  ( .a(\r125/LTV1 [41]), .b(\r125/LTV2 [41]), .out(
        \r125/LTV [42]) );
  xor2 \r125/UEQI_42  ( .a(N176), .b(N112), .out(n2519) );
  nand2 \r125/UGTI0_42  ( .a(n2518), .b(N176), .out(\r125/GTV1 [42]) );
  nand2 \r125/UGTI1_42  ( .a(\r125/AEQB [42]), .b(\r125/GTV [42]), .out(
        \r125/GTV2 [42]) );
  nand2 \r125/UGTI2_42  ( .a(\r125/GTV1 [42]), .b(\r125/GTV2 [42]), .out(
        \r125/GTV [43]) );
  nand2 \r125/ULTI0_42  ( .a(n2517), .b(N112), .out(\r125/LTV1 [42]) );
  nand2 \r125/ULTI1_42  ( .a(\r125/AEQB [42]), .b(\r125/LTV [42]), .out(
        \r125/LTV2 [42]) );
  nand2 \r125/ULTI2_42  ( .a(\r125/LTV1 [42]), .b(\r125/LTV2 [42]), .out(
        \r125/LTV [43]) );
  xor2 \r125/UEQI_43  ( .a(N175), .b(N111), .out(n2516) );
  nand2 \r125/UGTI0_43  ( .a(n2515), .b(N175), .out(\r125/GTV1 [43]) );
  nand2 \r125/UGTI1_43  ( .a(\r125/AEQB [43]), .b(\r125/GTV [43]), .out(
        \r125/GTV2 [43]) );
  nand2 \r125/UGTI2_43  ( .a(\r125/GTV1 [43]), .b(\r125/GTV2 [43]), .out(
        \r125/GTV [44]) );
  nand2 \r125/ULTI0_43  ( .a(n2514), .b(N111), .out(\r125/LTV1 [43]) );
  nand2 \r125/ULTI1_43  ( .a(\r125/AEQB [43]), .b(\r125/LTV [43]), .out(
        \r125/LTV2 [43]) );
  nand2 \r125/ULTI2_43  ( .a(\r125/LTV1 [43]), .b(\r125/LTV2 [43]), .out(
        \r125/LTV [44]) );
  xor2 \r125/UEQI_44  ( .a(N174), .b(N110), .out(n2513) );
  nand2 \r125/UGTI0_44  ( .a(n2512), .b(N174), .out(\r125/GTV1 [44]) );
  nand2 \r125/UGTI1_44  ( .a(\r125/AEQB [44]), .b(\r125/GTV [44]), .out(
        \r125/GTV2 [44]) );
  nand2 \r125/UGTI2_44  ( .a(\r125/GTV1 [44]), .b(\r125/GTV2 [44]), .out(
        \r125/GTV [45]) );
  nand2 \r125/ULTI0_44  ( .a(n2511), .b(N110), .out(\r125/LTV1 [44]) );
  nand2 \r125/ULTI1_44  ( .a(\r125/AEQB [44]), .b(\r125/LTV [44]), .out(
        \r125/LTV2 [44]) );
  nand2 \r125/ULTI2_44  ( .a(\r125/LTV1 [44]), .b(\r125/LTV2 [44]), .out(
        \r125/LTV [45]) );
  xor2 \r125/UEQI_45  ( .a(N173), .b(N109), .out(n2510) );
  nand2 \r125/UGTI0_45  ( .a(n2509), .b(N173), .out(\r125/GTV1 [45]) );
  nand2 \r125/UGTI1_45  ( .a(\r125/AEQB [45]), .b(\r125/GTV [45]), .out(
        \r125/GTV2 [45]) );
  nand2 \r125/UGTI2_45  ( .a(\r125/GTV1 [45]), .b(\r125/GTV2 [45]), .out(
        \r125/GTV [46]) );
  nand2 \r125/ULTI0_45  ( .a(n2508), .b(N109), .out(\r125/LTV1 [45]) );
  nand2 \r125/ULTI1_45  ( .a(\r125/AEQB [45]), .b(\r125/LTV [45]), .out(
        \r125/LTV2 [45]) );
  nand2 \r125/ULTI2_45  ( .a(\r125/LTV1 [45]), .b(\r125/LTV2 [45]), .out(
        \r125/LTV [46]) );
  xor2 \r125/UEQI_46  ( .a(N172), .b(N108), .out(n2507) );
  nand2 \r125/UGTI0_46  ( .a(n2506), .b(N172), .out(\r125/GTV1 [46]) );
  nand2 \r125/UGTI1_46  ( .a(\r125/AEQB [46]), .b(\r125/GTV [46]), .out(
        \r125/GTV2 [46]) );
  nand2 \r125/UGTI2_46  ( .a(\r125/GTV1 [46]), .b(\r125/GTV2 [46]), .out(
        \r125/GTV [47]) );
  nand2 \r125/ULTI0_46  ( .a(n2505), .b(N108), .out(\r125/LTV1 [46]) );
  nand2 \r125/ULTI1_46  ( .a(\r125/AEQB [46]), .b(\r125/LTV [46]), .out(
        \r125/LTV2 [46]) );
  nand2 \r125/ULTI2_46  ( .a(\r125/LTV1 [46]), .b(\r125/LTV2 [46]), .out(
        \r125/LTV [47]) );
  xor2 \r125/UEQI_47  ( .a(N171), .b(N107), .out(n2504) );
  nand2 \r125/UGTI0_47  ( .a(n2503), .b(N171), .out(\r125/GTV1 [47]) );
  nand2 \r125/UGTI1_47  ( .a(\r125/AEQB [47]), .b(\r125/GTV [47]), .out(
        \r125/GTV2 [47]) );
  nand2 \r125/UGTI2_47  ( .a(\r125/GTV1 [47]), .b(\r125/GTV2 [47]), .out(
        \r125/GTV [48]) );
  nand2 \r125/ULTI0_47  ( .a(n2502), .b(N107), .out(\r125/LTV1 [47]) );
  nand2 \r125/ULTI1_47  ( .a(\r125/AEQB [47]), .b(\r125/LTV [47]), .out(
        \r125/LTV2 [47]) );
  nand2 \r125/ULTI2_47  ( .a(\r125/LTV1 [47]), .b(\r125/LTV2 [47]), .out(
        \r125/LTV [48]) );
  xor2 \r125/UEQI_48  ( .a(N170), .b(N106), .out(n2501) );
  nand2 \r125/UGTI0_48  ( .a(n2500), .b(N170), .out(\r125/GTV1 [48]) );
  nand2 \r125/UGTI1_48  ( .a(\r125/AEQB [48]), .b(\r125/GTV [48]), .out(
        \r125/GTV2 [48]) );
  nand2 \r125/UGTI2_48  ( .a(\r125/GTV1 [48]), .b(\r125/GTV2 [48]), .out(
        \r125/GTV [49]) );
  nand2 \r125/ULTI0_48  ( .a(n2499), .b(N106), .out(\r125/LTV1 [48]) );
  nand2 \r125/ULTI1_48  ( .a(\r125/AEQB [48]), .b(\r125/LTV [48]), .out(
        \r125/LTV2 [48]) );
  nand2 \r125/ULTI2_48  ( .a(\r125/LTV1 [48]), .b(\r125/LTV2 [48]), .out(
        \r125/LTV [49]) );
  xor2 \r125/UEQI_49  ( .a(N169), .b(N105), .out(n2498) );
  nand2 \r125/UGTI0_49  ( .a(n2497), .b(N169), .out(\r125/GTV1 [49]) );
  nand2 \r125/UGTI1_49  ( .a(\r125/AEQB [49]), .b(\r125/GTV [49]), .out(
        \r125/GTV2 [49]) );
  nand2 \r125/UGTI2_49  ( .a(\r125/GTV1 [49]), .b(\r125/GTV2 [49]), .out(
        \r125/GTV [50]) );
  nand2 \r125/ULTI0_49  ( .a(n2496), .b(N105), .out(\r125/LTV1 [49]) );
  nand2 \r125/ULTI1_49  ( .a(\r125/AEQB [49]), .b(\r125/LTV [49]), .out(
        \r125/LTV2 [49]) );
  nand2 \r125/ULTI2_49  ( .a(\r125/LTV1 [49]), .b(\r125/LTV2 [49]), .out(
        \r125/LTV [50]) );
  xor2 \r125/UEQI_50  ( .a(N168), .b(N104), .out(n2495) );
  nand2 \r125/UGTI0_50  ( .a(n2494), .b(N168), .out(\r125/GTV1 [50]) );
  nand2 \r125/UGTI1_50  ( .a(\r125/AEQB [50]), .b(\r125/GTV [50]), .out(
        \r125/GTV2 [50]) );
  nand2 \r125/UGTI2_50  ( .a(\r125/GTV1 [50]), .b(\r125/GTV2 [50]), .out(
        \r125/GTV [51]) );
  nand2 \r125/ULTI0_50  ( .a(n2493), .b(N104), .out(\r125/LTV1 [50]) );
  nand2 \r125/ULTI1_50  ( .a(\r125/AEQB [50]), .b(\r125/LTV [50]), .out(
        \r125/LTV2 [50]) );
  nand2 \r125/ULTI2_50  ( .a(\r125/LTV1 [50]), .b(\r125/LTV2 [50]), .out(
        \r125/LTV [51]) );
  xor2 \r125/UEQI_51  ( .a(N167), .b(N103), .out(n2492) );
  nand2 \r125/UGTI0_51  ( .a(n2491), .b(N167), .out(\r125/GTV1 [51]) );
  nand2 \r125/UGTI1_51  ( .a(\r125/AEQB [51]), .b(\r125/GTV [51]), .out(
        \r125/GTV2 [51]) );
  nand2 \r125/UGTI2_51  ( .a(\r125/GTV1 [51]), .b(\r125/GTV2 [51]), .out(
        \r125/GTV [52]) );
  nand2 \r125/ULTI0_51  ( .a(n2490), .b(N103), .out(\r125/LTV1 [51]) );
  nand2 \r125/ULTI1_51  ( .a(\r125/AEQB [51]), .b(\r125/LTV [51]), .out(
        \r125/LTV2 [51]) );
  nand2 \r125/ULTI2_51  ( .a(\r125/LTV1 [51]), .b(\r125/LTV2 [51]), .out(
        \r125/LTV [52]) );
  xor2 \r125/UEQI_52  ( .a(N166), .b(N102), .out(n2489) );
  nand2 \r125/UGTI0_52  ( .a(n2488), .b(N166), .out(\r125/GTV1 [52]) );
  nand2 \r125/UGTI1_52  ( .a(\r125/AEQB [52]), .b(\r125/GTV [52]), .out(
        \r125/GTV2 [52]) );
  nand2 \r125/UGTI2_52  ( .a(\r125/GTV1 [52]), .b(\r125/GTV2 [52]), .out(
        \r125/GTV [53]) );
  nand2 \r125/ULTI0_52  ( .a(n2487), .b(N102), .out(\r125/LTV1 [52]) );
  nand2 \r125/ULTI1_52  ( .a(\r125/AEQB [52]), .b(\r125/LTV [52]), .out(
        \r125/LTV2 [52]) );
  nand2 \r125/ULTI2_52  ( .a(\r125/LTV1 [52]), .b(\r125/LTV2 [52]), .out(
        \r125/LTV [53]) );
  xor2 \r125/UEQI_53  ( .a(N165), .b(N101), .out(n2486) );
  nand2 \r125/UGTI0_53  ( .a(n2485), .b(N165), .out(\r125/GTV1 [53]) );
  nand2 \r125/UGTI1_53  ( .a(\r125/AEQB [53]), .b(\r125/GTV [53]), .out(
        \r125/GTV2 [53]) );
  nand2 \r125/UGTI2_53  ( .a(\r125/GTV1 [53]), .b(\r125/GTV2 [53]), .out(
        \r125/GTV [54]) );
  nand2 \r125/ULTI0_53  ( .a(n2484), .b(N101), .out(\r125/LTV1 [53]) );
  nand2 \r125/ULTI1_53  ( .a(\r125/AEQB [53]), .b(\r125/LTV [53]), .out(
        \r125/LTV2 [53]) );
  nand2 \r125/ULTI2_53  ( .a(\r125/LTV1 [53]), .b(\r125/LTV2 [53]), .out(
        \r125/LTV [54]) );
  xor2 \r125/UEQI_54  ( .a(N164), .b(N100), .out(n2483) );
  nand2 \r125/UGTI0_54  ( .a(n2482), .b(N164), .out(\r125/GTV1 [54]) );
  nand2 \r125/UGTI1_54  ( .a(\r125/AEQB [54]), .b(\r125/GTV [54]), .out(
        \r125/GTV2 [54]) );
  nand2 \r125/UGTI2_54  ( .a(\r125/GTV1 [54]), .b(\r125/GTV2 [54]), .out(
        \r125/GTV [55]) );
  nand2 \r125/ULTI0_54  ( .a(n2481), .b(N100), .out(\r125/LTV1 [54]) );
  nand2 \r125/ULTI1_54  ( .a(\r125/AEQB [54]), .b(\r125/LTV [54]), .out(
        \r125/LTV2 [54]) );
  nand2 \r125/ULTI2_54  ( .a(\r125/LTV1 [54]), .b(\r125/LTV2 [54]), .out(
        \r125/LTV [55]) );
  xor2 \r125/UEQI_55  ( .a(N163), .b(N99), .out(n2480) );
  nand2 \r125/UGTI0_55  ( .a(n2479), .b(N163), .out(\r125/GTV1 [55]) );
  nand2 \r125/UGTI1_55  ( .a(\r125/AEQB [55]), .b(\r125/GTV [55]), .out(
        \r125/GTV2 [55]) );
  nand2 \r125/UGTI2_55  ( .a(\r125/GTV1 [55]), .b(\r125/GTV2 [55]), .out(
        \r125/GTV [56]) );
  nand2 \r125/ULTI0_55  ( .a(n2478), .b(N99), .out(\r125/LTV1 [55]) );
  nand2 \r125/ULTI1_55  ( .a(\r125/AEQB [55]), .b(\r125/LTV [55]), .out(
        \r125/LTV2 [55]) );
  nand2 \r125/ULTI2_55  ( .a(\r125/LTV1 [55]), .b(\r125/LTV2 [55]), .out(
        \r125/LTV [56]) );
  xor2 \r125/UEQI_56  ( .a(N162), .b(N98), .out(n2477) );
  nand2 \r125/UGTI0_56  ( .a(n2476), .b(N162), .out(\r125/GTV1 [56]) );
  nand2 \r125/UGTI1_56  ( .a(\r125/AEQB [56]), .b(\r125/GTV [56]), .out(
        \r125/GTV2 [56]) );
  nand2 \r125/UGTI2_56  ( .a(\r125/GTV1 [56]), .b(\r125/GTV2 [56]), .out(
        \r125/GTV [57]) );
  nand2 \r125/ULTI0_56  ( .a(n2475), .b(N98), .out(\r125/LTV1 [56]) );
  nand2 \r125/ULTI1_56  ( .a(\r125/AEQB [56]), .b(\r125/LTV [56]), .out(
        \r125/LTV2 [56]) );
  nand2 \r125/ULTI2_56  ( .a(\r125/LTV1 [56]), .b(\r125/LTV2 [56]), .out(
        \r125/LTV [57]) );
  xor2 \r125/UEQI_57  ( .a(N161), .b(N97), .out(n2474) );
  nand2 \r125/UGTI0_57  ( .a(n2473), .b(N161), .out(\r125/GTV1 [57]) );
  nand2 \r125/UGTI1_57  ( .a(\r125/AEQB [57]), .b(\r125/GTV [57]), .out(
        \r125/GTV2 [57]) );
  nand2 \r125/UGTI2_57  ( .a(\r125/GTV1 [57]), .b(\r125/GTV2 [57]), .out(
        \r125/GTV [58]) );
  nand2 \r125/ULTI0_57  ( .a(n2472), .b(N97), .out(\r125/LTV1 [57]) );
  nand2 \r125/ULTI1_57  ( .a(\r125/AEQB [57]), .b(\r125/LTV [57]), .out(
        \r125/LTV2 [57]) );
  nand2 \r125/ULTI2_57  ( .a(\r125/LTV1 [57]), .b(\r125/LTV2 [57]), .out(
        \r125/LTV [58]) );
  xor2 \r125/UEQI_58  ( .a(N160), .b(N96), .out(n2471) );
  nand2 \r125/UGTI0_58  ( .a(n2470), .b(N160), .out(\r125/GTV1 [58]) );
  nand2 \r125/UGTI1_58  ( .a(\r125/AEQB [58]), .b(\r125/GTV [58]), .out(
        \r125/GTV2 [58]) );
  nand2 \r125/UGTI2_58  ( .a(\r125/GTV1 [58]), .b(\r125/GTV2 [58]), .out(
        \r125/GTV [59]) );
  nand2 \r125/ULTI0_58  ( .a(n2469), .b(N96), .out(\r125/LTV1 [58]) );
  nand2 \r125/ULTI1_58  ( .a(\r125/AEQB [58]), .b(\r125/LTV [58]), .out(
        \r125/LTV2 [58]) );
  nand2 \r125/ULTI2_58  ( .a(\r125/LTV1 [58]), .b(\r125/LTV2 [58]), .out(
        \r125/LTV [59]) );
  xor2 \r125/UEQI_59  ( .a(N159), .b(N95), .out(n2468) );
  nand2 \r125/UGTI0_59  ( .a(n2467), .b(N159), .out(\r125/GTV1 [59]) );
  nand2 \r125/UGTI1_59  ( .a(\r125/AEQB [59]), .b(\r125/GTV [59]), .out(
        \r125/GTV2 [59]) );
  nand2 \r125/UGTI2_59  ( .a(\r125/GTV1 [59]), .b(\r125/GTV2 [59]), .out(
        \r125/GTV [60]) );
  nand2 \r125/ULTI0_59  ( .a(n2466), .b(N95), .out(\r125/LTV1 [59]) );
  nand2 \r125/ULTI1_59  ( .a(\r125/AEQB [59]), .b(\r125/LTV [59]), .out(
        \r125/LTV2 [59]) );
  nand2 \r125/ULTI2_59  ( .a(\r125/LTV1 [59]), .b(\r125/LTV2 [59]), .out(
        \r125/LTV [60]) );
  xor2 \r125/UEQI_60  ( .a(N158), .b(N94), .out(n2465) );
  nand2 \r125/UGTI0_60  ( .a(n2464), .b(N158), .out(\r125/GTV1 [60]) );
  nand2 \r125/UGTI1_60  ( .a(\r125/AEQB [60]), .b(\r125/GTV [60]), .out(
        \r125/GTV2 [60]) );
  nand2 \r125/UGTI2_60  ( .a(\r125/GTV1 [60]), .b(\r125/GTV2 [60]), .out(
        \r125/GTV [61]) );
  nand2 \r125/ULTI0_60  ( .a(n2463), .b(N94), .out(\r125/LTV1 [60]) );
  nand2 \r125/ULTI1_60  ( .a(\r125/AEQB [60]), .b(\r125/LTV [60]), .out(
        \r125/LTV2 [60]) );
  nand2 \r125/ULTI2_60  ( .a(\r125/LTV1 [60]), .b(\r125/LTV2 [60]), .out(
        \r125/LTV [61]) );
  xor2 \r125/UEQI_61  ( .a(N157), .b(N93), .out(n2462) );
  nand2 \r125/UGTI0_61  ( .a(n2461), .b(N157), .out(\r125/GTV1 [61]) );
  nand2 \r125/UGTI1_61  ( .a(\r125/AEQB [61]), .b(\r125/GTV [61]), .out(
        \r125/GTV2 [61]) );
  nand2 \r125/UGTI2_61  ( .a(\r125/GTV1 [61]), .b(\r125/GTV2 [61]), .out(
        \r125/GTV [62]) );
  nand2 \r125/ULTI0_61  ( .a(n2460), .b(N93), .out(\r125/LTV1 [61]) );
  nand2 \r125/ULTI1_61  ( .a(\r125/AEQB [61]), .b(\r125/LTV [61]), .out(
        \r125/LTV2 [61]) );
  nand2 \r125/ULTI2_61  ( .a(\r125/LTV1 [61]), .b(\r125/LTV2 [61]), .out(
        \r125/LTV [62]) );
  xor2 \r125/UEQI_62  ( .a(N156), .b(N92), .out(n2459) );
  nand2 \r125/UGTI0_62  ( .a(n2458), .b(N156), .out(\r125/GTV1 [62]) );
  nand2 \r125/UGTI1_62  ( .a(\r125/AEQB [62]), .b(\r125/GTV [62]), .out(
        \r125/GTV2 [62]) );
  nand2 \r125/UGTI2_62  ( .a(\r125/GTV1 [62]), .b(\r125/GTV2 [62]), .out(
        \r125/GTV [63]) );
  nand2 \r125/ULTI0_62  ( .a(n2457), .b(N92), .out(\r125/LTV1 [62]) );
  nand2 \r125/ULTI1_62  ( .a(\r125/AEQB [62]), .b(\r125/LTV [62]), .out(
        \r125/LTV2 [62]) );
  nand2 \r125/ULTI2_62  ( .a(\r125/LTV1 [62]), .b(\r125/LTV2 [62]), .out(
        \r125/LTV [63]) );
  nor2 \eq_47_3/UEQ  ( .a(\eq_47_3/GT ), .b(\eq_47_3/LT ), .out(N16) );
  nand2 \eq_47_3/UNGT0  ( .a(current_floor_output_elevator2[0]), .b(n2456), 
        .out(n2455) );
  nand2 \eq_47_3/UNLT0  ( .a(destination_floor_elevator2[0]), .b(n2454), .out(
        n2453) );
  xor2 \eq_47_3/UEQI  ( .a(\eq_47_3/SA ), .b(\eq_47_3/SB ), .out(n2452) );
  nand2 \eq_47_3/UGTI0  ( .a(n2451), .b(\eq_47_3/SA ), .out(\eq_47_3/GTV1 [63]) );
  nand2 \eq_47_3/UGTI1  ( .a(\eq_47_3/AEQB [63]), .b(\eq_47_3/GTV [63]), .out(
        \eq_47_3/GTV2 [63]) );
  nand2 \eq_47_3/UGTI2  ( .a(\eq_47_3/GTV1 [63]), .b(\eq_47_3/GTV2 [63]), 
        .out(\eq_47_3/GT ) );
  nand2 \eq_47_3/ULTI0  ( .a(n2450), .b(\eq_47_3/SB ), .out(\eq_47_3/LTV1 [63]) );
  nand2 \eq_47_3/ULTI1  ( .a(\eq_47_3/AEQB [63]), .b(\eq_47_3/LTV [63]), .out(
        \eq_47_3/LTV2 [63]) );
  nand2 \eq_47_3/ULTI2  ( .a(\eq_47_3/LTV1 [63]), .b(\eq_47_3/LTV2 [63]), 
        .out(\eq_47_3/LT ) );
  xor2 \eq_47_3/UEQI_1  ( .a(current_floor_output_elevator2[1]), .b(
        destination_floor_elevator2[1]), .out(n2449) );
  nand2 \eq_47_3/UGTI0_1  ( .a(n2448), .b(current_floor_output_elevator2[1]), 
        .out(\eq_47_3/GTV1 [1]) );
  nand2 \eq_47_3/UGTI1_1  ( .a(\eq_47_3/AEQB [1]), .b(\eq_47_3/GTV [1]), .out(
        \eq_47_3/GTV2 [1]) );
  nand2 \eq_47_3/UGTI2_1  ( .a(\eq_47_3/GTV1 [1]), .b(\eq_47_3/GTV2 [1]), 
        .out(\eq_47_3/GTV [2]) );
  nand2 \eq_47_3/ULTI0_1  ( .a(n2447), .b(destination_floor_elevator2[1]), 
        .out(\eq_47_3/LTV1 [1]) );
  nand2 \eq_47_3/ULTI1_1  ( .a(\eq_47_3/AEQB [1]), .b(\eq_47_3/LTV [1]), .out(
        \eq_47_3/LTV2 [1]) );
  nand2 \eq_47_3/ULTI2_1  ( .a(\eq_47_3/LTV1 [1]), .b(\eq_47_3/LTV2 [1]), 
        .out(\eq_47_3/LTV [2]) );
  xor2 \eq_47_3/UEQI_2  ( .a(current_floor_output_elevator2[2]), .b(
        destination_floor_elevator2[2]), .out(n2446) );
  nand2 \eq_47_3/UGTI0_2  ( .a(n2445), .b(current_floor_output_elevator2[2]), 
        .out(\eq_47_3/GTV1 [2]) );
  nand2 \eq_47_3/UGTI1_2  ( .a(\eq_47_3/AEQB [2]), .b(\eq_47_3/GTV [2]), .out(
        \eq_47_3/GTV2 [2]) );
  nand2 \eq_47_3/UGTI2_2  ( .a(\eq_47_3/GTV1 [2]), .b(\eq_47_3/GTV2 [2]), 
        .out(\eq_47_3/GTV [3]) );
  nand2 \eq_47_3/ULTI0_2  ( .a(n2444), .b(destination_floor_elevator2[2]), 
        .out(\eq_47_3/LTV1 [2]) );
  nand2 \eq_47_3/ULTI1_2  ( .a(\eq_47_3/AEQB [2]), .b(\eq_47_3/LTV [2]), .out(
        \eq_47_3/LTV2 [2]) );
  nand2 \eq_47_3/ULTI2_2  ( .a(\eq_47_3/LTV1 [2]), .b(\eq_47_3/LTV2 [2]), 
        .out(\eq_47_3/LTV [3]) );
  xor2 \eq_47_3/UEQI_3  ( .a(current_floor_output_elevator2[3]), .b(
        destination_floor_elevator2[3]), .out(n2443) );
  nand2 \eq_47_3/UGTI0_3  ( .a(n2442), .b(current_floor_output_elevator2[3]), 
        .out(\eq_47_3/GTV1 [3]) );
  nand2 \eq_47_3/UGTI1_3  ( .a(\eq_47_3/AEQB [3]), .b(\eq_47_3/GTV [3]), .out(
        \eq_47_3/GTV2 [3]) );
  nand2 \eq_47_3/UGTI2_3  ( .a(\eq_47_3/GTV1 [3]), .b(\eq_47_3/GTV2 [3]), 
        .out(\eq_47_3/GTV [4]) );
  nand2 \eq_47_3/ULTI0_3  ( .a(n2441), .b(destination_floor_elevator2[3]), 
        .out(\eq_47_3/LTV1 [3]) );
  nand2 \eq_47_3/ULTI1_3  ( .a(\eq_47_3/AEQB [3]), .b(\eq_47_3/LTV [3]), .out(
        \eq_47_3/LTV2 [3]) );
  nand2 \eq_47_3/ULTI2_3  ( .a(\eq_47_3/LTV1 [3]), .b(\eq_47_3/LTV2 [3]), 
        .out(\eq_47_3/LTV [4]) );
  xor2 \eq_47_3/UEQI_4  ( .a(current_floor_output_elevator2[4]), .b(
        destination_floor_elevator2[4]), .out(n2440) );
  nand2 \eq_47_3/UGTI0_4  ( .a(n2439), .b(current_floor_output_elevator2[4]), 
        .out(\eq_47_3/GTV1 [4]) );
  nand2 \eq_47_3/UGTI1_4  ( .a(\eq_47_3/AEQB [4]), .b(\eq_47_3/GTV [4]), .out(
        \eq_47_3/GTV2 [4]) );
  nand2 \eq_47_3/UGTI2_4  ( .a(\eq_47_3/GTV1 [4]), .b(\eq_47_3/GTV2 [4]), 
        .out(\eq_47_3/GTV [5]) );
  nand2 \eq_47_3/ULTI0_4  ( .a(n2438), .b(destination_floor_elevator2[4]), 
        .out(\eq_47_3/LTV1 [4]) );
  nand2 \eq_47_3/ULTI1_4  ( .a(\eq_47_3/AEQB [4]), .b(\eq_47_3/LTV [4]), .out(
        \eq_47_3/LTV2 [4]) );
  nand2 \eq_47_3/ULTI2_4  ( .a(\eq_47_3/LTV1 [4]), .b(\eq_47_3/LTV2 [4]), 
        .out(\eq_47_3/LTV [5]) );
  xor2 \eq_47_3/UEQI_5  ( .a(current_floor_output_elevator2[5]), .b(
        destination_floor_elevator2[5]), .out(n2437) );
  nand2 \eq_47_3/UGTI0_5  ( .a(n2436), .b(current_floor_output_elevator2[5]), 
        .out(\eq_47_3/GTV1 [5]) );
  nand2 \eq_47_3/UGTI1_5  ( .a(\eq_47_3/AEQB [5]), .b(\eq_47_3/GTV [5]), .out(
        \eq_47_3/GTV2 [5]) );
  nand2 \eq_47_3/UGTI2_5  ( .a(\eq_47_3/GTV1 [5]), .b(\eq_47_3/GTV2 [5]), 
        .out(\eq_47_3/GTV [6]) );
  nand2 \eq_47_3/ULTI0_5  ( .a(n2435), .b(destination_floor_elevator2[5]), 
        .out(\eq_47_3/LTV1 [5]) );
  nand2 \eq_47_3/ULTI1_5  ( .a(\eq_47_3/AEQB [5]), .b(\eq_47_3/LTV [5]), .out(
        \eq_47_3/LTV2 [5]) );
  nand2 \eq_47_3/ULTI2_5  ( .a(\eq_47_3/LTV1 [5]), .b(\eq_47_3/LTV2 [5]), 
        .out(\eq_47_3/LTV [6]) );
  xor2 \eq_47_3/UEQI_6  ( .a(current_floor_output_elevator2[6]), .b(
        destination_floor_elevator2[6]), .out(n2434) );
  nand2 \eq_47_3/UGTI0_6  ( .a(n2433), .b(current_floor_output_elevator2[6]), 
        .out(\eq_47_3/GTV1 [6]) );
  nand2 \eq_47_3/UGTI1_6  ( .a(\eq_47_3/AEQB [6]), .b(\eq_47_3/GTV [6]), .out(
        \eq_47_3/GTV2 [6]) );
  nand2 \eq_47_3/UGTI2_6  ( .a(\eq_47_3/GTV1 [6]), .b(\eq_47_3/GTV2 [6]), 
        .out(\eq_47_3/GTV [7]) );
  nand2 \eq_47_3/ULTI0_6  ( .a(n2432), .b(destination_floor_elevator2[6]), 
        .out(\eq_47_3/LTV1 [6]) );
  nand2 \eq_47_3/ULTI1_6  ( .a(\eq_47_3/AEQB [6]), .b(\eq_47_3/LTV [6]), .out(
        \eq_47_3/LTV2 [6]) );
  nand2 \eq_47_3/ULTI2_6  ( .a(\eq_47_3/LTV1 [6]), .b(\eq_47_3/LTV2 [6]), 
        .out(\eq_47_3/LTV [7]) );
  xor2 \eq_47_3/UEQI_7  ( .a(current_floor_output_elevator2[7]), .b(
        destination_floor_elevator2[7]), .out(n2431) );
  nand2 \eq_47_3/UGTI0_7  ( .a(n2430), .b(current_floor_output_elevator2[7]), 
        .out(\eq_47_3/GTV1 [7]) );
  nand2 \eq_47_3/UGTI1_7  ( .a(\eq_47_3/AEQB [7]), .b(\eq_47_3/GTV [7]), .out(
        \eq_47_3/GTV2 [7]) );
  nand2 \eq_47_3/UGTI2_7  ( .a(\eq_47_3/GTV1 [7]), .b(\eq_47_3/GTV2 [7]), 
        .out(\eq_47_3/GTV [8]) );
  nand2 \eq_47_3/ULTI0_7  ( .a(n2429), .b(destination_floor_elevator2[7]), 
        .out(\eq_47_3/LTV1 [7]) );
  nand2 \eq_47_3/ULTI1_7  ( .a(\eq_47_3/AEQB [7]), .b(\eq_47_3/LTV [7]), .out(
        \eq_47_3/LTV2 [7]) );
  nand2 \eq_47_3/ULTI2_7  ( .a(\eq_47_3/LTV1 [7]), .b(\eq_47_3/LTV2 [7]), 
        .out(\eq_47_3/LTV [8]) );
  xor2 \eq_47_3/UEQI_8  ( .a(current_floor_output_elevator2[8]), .b(
        destination_floor_elevator2[8]), .out(n2428) );
  nand2 \eq_47_3/UGTI0_8  ( .a(n2427), .b(current_floor_output_elevator2[8]), 
        .out(\eq_47_3/GTV1 [8]) );
  nand2 \eq_47_3/UGTI1_8  ( .a(\eq_47_3/AEQB [8]), .b(\eq_47_3/GTV [8]), .out(
        \eq_47_3/GTV2 [8]) );
  nand2 \eq_47_3/UGTI2_8  ( .a(\eq_47_3/GTV1 [8]), .b(\eq_47_3/GTV2 [8]), 
        .out(\eq_47_3/GTV [9]) );
  nand2 \eq_47_3/ULTI0_8  ( .a(n2426), .b(destination_floor_elevator2[8]), 
        .out(\eq_47_3/LTV1 [8]) );
  nand2 \eq_47_3/ULTI1_8  ( .a(\eq_47_3/AEQB [8]), .b(\eq_47_3/LTV [8]), .out(
        \eq_47_3/LTV2 [8]) );
  nand2 \eq_47_3/ULTI2_8  ( .a(\eq_47_3/LTV1 [8]), .b(\eq_47_3/LTV2 [8]), 
        .out(\eq_47_3/LTV [9]) );
  xor2 \eq_47_3/UEQI_9  ( .a(current_floor_output_elevator2[9]), .b(
        destination_floor_elevator2[9]), .out(n2425) );
  nand2 \eq_47_3/UGTI0_9  ( .a(n2424), .b(current_floor_output_elevator2[9]), 
        .out(\eq_47_3/GTV1 [9]) );
  nand2 \eq_47_3/UGTI1_9  ( .a(\eq_47_3/AEQB [9]), .b(\eq_47_3/GTV [9]), .out(
        \eq_47_3/GTV2 [9]) );
  nand2 \eq_47_3/UGTI2_9  ( .a(\eq_47_3/GTV1 [9]), .b(\eq_47_3/GTV2 [9]), 
        .out(\eq_47_3/GTV [10]) );
  nand2 \eq_47_3/ULTI0_9  ( .a(n2423), .b(destination_floor_elevator2[9]), 
        .out(\eq_47_3/LTV1 [9]) );
  nand2 \eq_47_3/ULTI1_9  ( .a(\eq_47_3/AEQB [9]), .b(\eq_47_3/LTV [9]), .out(
        \eq_47_3/LTV2 [9]) );
  nand2 \eq_47_3/ULTI2_9  ( .a(\eq_47_3/LTV1 [9]), .b(\eq_47_3/LTV2 [9]), 
        .out(\eq_47_3/LTV [10]) );
  xor2 \eq_47_3/UEQI_10  ( .a(current_floor_output_elevator2[10]), .b(
        destination_floor_elevator2[10]), .out(n2422) );
  nand2 \eq_47_3/UGTI0_10  ( .a(n2421), .b(current_floor_output_elevator2[10]), 
        .out(\eq_47_3/GTV1 [10]) );
  nand2 \eq_47_3/UGTI1_10  ( .a(\eq_47_3/AEQB [10]), .b(\eq_47_3/GTV [10]), 
        .out(\eq_47_3/GTV2 [10]) );
  nand2 \eq_47_3/UGTI2_10  ( .a(\eq_47_3/GTV1 [10]), .b(\eq_47_3/GTV2 [10]), 
        .out(\eq_47_3/GTV [11]) );
  nand2 \eq_47_3/ULTI0_10  ( .a(n2420), .b(destination_floor_elevator2[10]), 
        .out(\eq_47_3/LTV1 [10]) );
  nand2 \eq_47_3/ULTI1_10  ( .a(\eq_47_3/AEQB [10]), .b(\eq_47_3/LTV [10]), 
        .out(\eq_47_3/LTV2 [10]) );
  nand2 \eq_47_3/ULTI2_10  ( .a(\eq_47_3/LTV1 [10]), .b(\eq_47_3/LTV2 [10]), 
        .out(\eq_47_3/LTV [11]) );
  xor2 \eq_47_3/UEQI_11  ( .a(current_floor_output_elevator2[11]), .b(
        destination_floor_elevator2[11]), .out(n2419) );
  nand2 \eq_47_3/UGTI0_11  ( .a(n2418), .b(current_floor_output_elevator2[11]), 
        .out(\eq_47_3/GTV1 [11]) );
  nand2 \eq_47_3/UGTI1_11  ( .a(\eq_47_3/AEQB [11]), .b(\eq_47_3/GTV [11]), 
        .out(\eq_47_3/GTV2 [11]) );
  nand2 \eq_47_3/UGTI2_11  ( .a(\eq_47_3/GTV1 [11]), .b(\eq_47_3/GTV2 [11]), 
        .out(\eq_47_3/GTV [12]) );
  nand2 \eq_47_3/ULTI0_11  ( .a(n2417), .b(destination_floor_elevator2[11]), 
        .out(\eq_47_3/LTV1 [11]) );
  nand2 \eq_47_3/ULTI1_11  ( .a(\eq_47_3/AEQB [11]), .b(\eq_47_3/LTV [11]), 
        .out(\eq_47_3/LTV2 [11]) );
  nand2 \eq_47_3/ULTI2_11  ( .a(\eq_47_3/LTV1 [11]), .b(\eq_47_3/LTV2 [11]), 
        .out(\eq_47_3/LTV [12]) );
  xor2 \eq_47_3/UEQI_12  ( .a(current_floor_output_elevator2[12]), .b(
        destination_floor_elevator2[12]), .out(n2416) );
  nand2 \eq_47_3/UGTI0_12  ( .a(n2415), .b(current_floor_output_elevator2[12]), 
        .out(\eq_47_3/GTV1 [12]) );
  nand2 \eq_47_3/UGTI1_12  ( .a(\eq_47_3/AEQB [12]), .b(\eq_47_3/GTV [12]), 
        .out(\eq_47_3/GTV2 [12]) );
  nand2 \eq_47_3/UGTI2_12  ( .a(\eq_47_3/GTV1 [12]), .b(\eq_47_3/GTV2 [12]), 
        .out(\eq_47_3/GTV [13]) );
  nand2 \eq_47_3/ULTI0_12  ( .a(n2414), .b(destination_floor_elevator2[12]), 
        .out(\eq_47_3/LTV1 [12]) );
  nand2 \eq_47_3/ULTI1_12  ( .a(\eq_47_3/AEQB [12]), .b(\eq_47_3/LTV [12]), 
        .out(\eq_47_3/LTV2 [12]) );
  nand2 \eq_47_3/ULTI2_12  ( .a(\eq_47_3/LTV1 [12]), .b(\eq_47_3/LTV2 [12]), 
        .out(\eq_47_3/LTV [13]) );
  xor2 \eq_47_3/UEQI_13  ( .a(current_floor_output_elevator2[13]), .b(
        destination_floor_elevator2[13]), .out(n2413) );
  nand2 \eq_47_3/UGTI0_13  ( .a(n2412), .b(current_floor_output_elevator2[13]), 
        .out(\eq_47_3/GTV1 [13]) );
  nand2 \eq_47_3/UGTI1_13  ( .a(\eq_47_3/AEQB [13]), .b(\eq_47_3/GTV [13]), 
        .out(\eq_47_3/GTV2 [13]) );
  nand2 \eq_47_3/UGTI2_13  ( .a(\eq_47_3/GTV1 [13]), .b(\eq_47_3/GTV2 [13]), 
        .out(\eq_47_3/GTV [14]) );
  nand2 \eq_47_3/ULTI0_13  ( .a(n2411), .b(destination_floor_elevator2[13]), 
        .out(\eq_47_3/LTV1 [13]) );
  nand2 \eq_47_3/ULTI1_13  ( .a(\eq_47_3/AEQB [13]), .b(\eq_47_3/LTV [13]), 
        .out(\eq_47_3/LTV2 [13]) );
  nand2 \eq_47_3/ULTI2_13  ( .a(\eq_47_3/LTV1 [13]), .b(\eq_47_3/LTV2 [13]), 
        .out(\eq_47_3/LTV [14]) );
  xor2 \eq_47_3/UEQI_14  ( .a(current_floor_output_elevator2[14]), .b(
        destination_floor_elevator2[14]), .out(n2410) );
  nand2 \eq_47_3/UGTI0_14  ( .a(n2409), .b(current_floor_output_elevator2[14]), 
        .out(\eq_47_3/GTV1 [14]) );
  nand2 \eq_47_3/UGTI1_14  ( .a(\eq_47_3/AEQB [14]), .b(\eq_47_3/GTV [14]), 
        .out(\eq_47_3/GTV2 [14]) );
  nand2 \eq_47_3/UGTI2_14  ( .a(\eq_47_3/GTV1 [14]), .b(\eq_47_3/GTV2 [14]), 
        .out(\eq_47_3/GTV [15]) );
  nand2 \eq_47_3/ULTI0_14  ( .a(n2408), .b(destination_floor_elevator2[14]), 
        .out(\eq_47_3/LTV1 [14]) );
  nand2 \eq_47_3/ULTI1_14  ( .a(\eq_47_3/AEQB [14]), .b(\eq_47_3/LTV [14]), 
        .out(\eq_47_3/LTV2 [14]) );
  nand2 \eq_47_3/ULTI2_14  ( .a(\eq_47_3/LTV1 [14]), .b(\eq_47_3/LTV2 [14]), 
        .out(\eq_47_3/LTV [15]) );
  xor2 \eq_47_3/UEQI_15  ( .a(current_floor_output_elevator2[15]), .b(
        destination_floor_elevator2[15]), .out(n2407) );
  nand2 \eq_47_3/UGTI0_15  ( .a(n2406), .b(current_floor_output_elevator2[15]), 
        .out(\eq_47_3/GTV1 [15]) );
  nand2 \eq_47_3/UGTI1_15  ( .a(\eq_47_3/AEQB [15]), .b(\eq_47_3/GTV [15]), 
        .out(\eq_47_3/GTV2 [15]) );
  nand2 \eq_47_3/UGTI2_15  ( .a(\eq_47_3/GTV1 [15]), .b(\eq_47_3/GTV2 [15]), 
        .out(\eq_47_3/GTV [16]) );
  nand2 \eq_47_3/ULTI0_15  ( .a(n2405), .b(destination_floor_elevator2[15]), 
        .out(\eq_47_3/LTV1 [15]) );
  nand2 \eq_47_3/ULTI1_15  ( .a(\eq_47_3/AEQB [15]), .b(\eq_47_3/LTV [15]), 
        .out(\eq_47_3/LTV2 [15]) );
  nand2 \eq_47_3/ULTI2_15  ( .a(\eq_47_3/LTV1 [15]), .b(\eq_47_3/LTV2 [15]), 
        .out(\eq_47_3/LTV [16]) );
  xor2 \eq_47_3/UEQI_16  ( .a(current_floor_output_elevator2[16]), .b(
        destination_floor_elevator2[16]), .out(n2404) );
  nand2 \eq_47_3/UGTI0_16  ( .a(n2403), .b(current_floor_output_elevator2[16]), 
        .out(\eq_47_3/GTV1 [16]) );
  nand2 \eq_47_3/UGTI1_16  ( .a(\eq_47_3/AEQB [16]), .b(\eq_47_3/GTV [16]), 
        .out(\eq_47_3/GTV2 [16]) );
  nand2 \eq_47_3/UGTI2_16  ( .a(\eq_47_3/GTV1 [16]), .b(\eq_47_3/GTV2 [16]), 
        .out(\eq_47_3/GTV [17]) );
  nand2 \eq_47_3/ULTI0_16  ( .a(n2402), .b(destination_floor_elevator2[16]), 
        .out(\eq_47_3/LTV1 [16]) );
  nand2 \eq_47_3/ULTI1_16  ( .a(\eq_47_3/AEQB [16]), .b(\eq_47_3/LTV [16]), 
        .out(\eq_47_3/LTV2 [16]) );
  nand2 \eq_47_3/ULTI2_16  ( .a(\eq_47_3/LTV1 [16]), .b(\eq_47_3/LTV2 [16]), 
        .out(\eq_47_3/LTV [17]) );
  xor2 \eq_47_3/UEQI_17  ( .a(current_floor_output_elevator2[17]), .b(
        destination_floor_elevator2[17]), .out(n2401) );
  nand2 \eq_47_3/UGTI0_17  ( .a(n2400), .b(current_floor_output_elevator2[17]), 
        .out(\eq_47_3/GTV1 [17]) );
  nand2 \eq_47_3/UGTI1_17  ( .a(\eq_47_3/AEQB [17]), .b(\eq_47_3/GTV [17]), 
        .out(\eq_47_3/GTV2 [17]) );
  nand2 \eq_47_3/UGTI2_17  ( .a(\eq_47_3/GTV1 [17]), .b(\eq_47_3/GTV2 [17]), 
        .out(\eq_47_3/GTV [18]) );
  nand2 \eq_47_3/ULTI0_17  ( .a(n2399), .b(destination_floor_elevator2[17]), 
        .out(\eq_47_3/LTV1 [17]) );
  nand2 \eq_47_3/ULTI1_17  ( .a(\eq_47_3/AEQB [17]), .b(\eq_47_3/LTV [17]), 
        .out(\eq_47_3/LTV2 [17]) );
  nand2 \eq_47_3/ULTI2_17  ( .a(\eq_47_3/LTV1 [17]), .b(\eq_47_3/LTV2 [17]), 
        .out(\eq_47_3/LTV [18]) );
  xor2 \eq_47_3/UEQI_18  ( .a(current_floor_output_elevator2[18]), .b(
        destination_floor_elevator2[18]), .out(n2398) );
  nand2 \eq_47_3/UGTI0_18  ( .a(n2397), .b(current_floor_output_elevator2[18]), 
        .out(\eq_47_3/GTV1 [18]) );
  nand2 \eq_47_3/UGTI1_18  ( .a(\eq_47_3/AEQB [18]), .b(\eq_47_3/GTV [18]), 
        .out(\eq_47_3/GTV2 [18]) );
  nand2 \eq_47_3/UGTI2_18  ( .a(\eq_47_3/GTV1 [18]), .b(\eq_47_3/GTV2 [18]), 
        .out(\eq_47_3/GTV [19]) );
  nand2 \eq_47_3/ULTI0_18  ( .a(n2396), .b(destination_floor_elevator2[18]), 
        .out(\eq_47_3/LTV1 [18]) );
  nand2 \eq_47_3/ULTI1_18  ( .a(\eq_47_3/AEQB [18]), .b(\eq_47_3/LTV [18]), 
        .out(\eq_47_3/LTV2 [18]) );
  nand2 \eq_47_3/ULTI2_18  ( .a(\eq_47_3/LTV1 [18]), .b(\eq_47_3/LTV2 [18]), 
        .out(\eq_47_3/LTV [19]) );
  xor2 \eq_47_3/UEQI_19  ( .a(current_floor_output_elevator2[19]), .b(
        destination_floor_elevator2[19]), .out(n2395) );
  nand2 \eq_47_3/UGTI0_19  ( .a(n2394), .b(current_floor_output_elevator2[19]), 
        .out(\eq_47_3/GTV1 [19]) );
  nand2 \eq_47_3/UGTI1_19  ( .a(\eq_47_3/AEQB [19]), .b(\eq_47_3/GTV [19]), 
        .out(\eq_47_3/GTV2 [19]) );
  nand2 \eq_47_3/UGTI2_19  ( .a(\eq_47_3/GTV1 [19]), .b(\eq_47_3/GTV2 [19]), 
        .out(\eq_47_3/GTV [20]) );
  nand2 \eq_47_3/ULTI0_19  ( .a(n2393), .b(destination_floor_elevator2[19]), 
        .out(\eq_47_3/LTV1 [19]) );
  nand2 \eq_47_3/ULTI1_19  ( .a(\eq_47_3/AEQB [19]), .b(\eq_47_3/LTV [19]), 
        .out(\eq_47_3/LTV2 [19]) );
  nand2 \eq_47_3/ULTI2_19  ( .a(\eq_47_3/LTV1 [19]), .b(\eq_47_3/LTV2 [19]), 
        .out(\eq_47_3/LTV [20]) );
  xor2 \eq_47_3/UEQI_20  ( .a(current_floor_output_elevator2[20]), .b(
        destination_floor_elevator2[20]), .out(n2392) );
  nand2 \eq_47_3/UGTI0_20  ( .a(n2391), .b(current_floor_output_elevator2[20]), 
        .out(\eq_47_3/GTV1 [20]) );
  nand2 \eq_47_3/UGTI1_20  ( .a(\eq_47_3/AEQB [20]), .b(\eq_47_3/GTV [20]), 
        .out(\eq_47_3/GTV2 [20]) );
  nand2 \eq_47_3/UGTI2_20  ( .a(\eq_47_3/GTV1 [20]), .b(\eq_47_3/GTV2 [20]), 
        .out(\eq_47_3/GTV [21]) );
  nand2 \eq_47_3/ULTI0_20  ( .a(n2390), .b(destination_floor_elevator2[20]), 
        .out(\eq_47_3/LTV1 [20]) );
  nand2 \eq_47_3/ULTI1_20  ( .a(\eq_47_3/AEQB [20]), .b(\eq_47_3/LTV [20]), 
        .out(\eq_47_3/LTV2 [20]) );
  nand2 \eq_47_3/ULTI2_20  ( .a(\eq_47_3/LTV1 [20]), .b(\eq_47_3/LTV2 [20]), 
        .out(\eq_47_3/LTV [21]) );
  xor2 \eq_47_3/UEQI_21  ( .a(current_floor_output_elevator2[21]), .b(
        destination_floor_elevator2[21]), .out(n2389) );
  nand2 \eq_47_3/UGTI0_21  ( .a(n2388), .b(current_floor_output_elevator2[21]), 
        .out(\eq_47_3/GTV1 [21]) );
  nand2 \eq_47_3/UGTI1_21  ( .a(\eq_47_3/AEQB [21]), .b(\eq_47_3/GTV [21]), 
        .out(\eq_47_3/GTV2 [21]) );
  nand2 \eq_47_3/UGTI2_21  ( .a(\eq_47_3/GTV1 [21]), .b(\eq_47_3/GTV2 [21]), 
        .out(\eq_47_3/GTV [22]) );
  nand2 \eq_47_3/ULTI0_21  ( .a(n2387), .b(destination_floor_elevator2[21]), 
        .out(\eq_47_3/LTV1 [21]) );
  nand2 \eq_47_3/ULTI1_21  ( .a(\eq_47_3/AEQB [21]), .b(\eq_47_3/LTV [21]), 
        .out(\eq_47_3/LTV2 [21]) );
  nand2 \eq_47_3/ULTI2_21  ( .a(\eq_47_3/LTV1 [21]), .b(\eq_47_3/LTV2 [21]), 
        .out(\eq_47_3/LTV [22]) );
  xor2 \eq_47_3/UEQI_22  ( .a(current_floor_output_elevator2[22]), .b(
        destination_floor_elevator2[22]), .out(n2386) );
  nand2 \eq_47_3/UGTI0_22  ( .a(n2385), .b(current_floor_output_elevator2[22]), 
        .out(\eq_47_3/GTV1 [22]) );
  nand2 \eq_47_3/UGTI1_22  ( .a(\eq_47_3/AEQB [22]), .b(\eq_47_3/GTV [22]), 
        .out(\eq_47_3/GTV2 [22]) );
  nand2 \eq_47_3/UGTI2_22  ( .a(\eq_47_3/GTV1 [22]), .b(\eq_47_3/GTV2 [22]), 
        .out(\eq_47_3/GTV [23]) );
  nand2 \eq_47_3/ULTI0_22  ( .a(n2384), .b(destination_floor_elevator2[22]), 
        .out(\eq_47_3/LTV1 [22]) );
  nand2 \eq_47_3/ULTI1_22  ( .a(\eq_47_3/AEQB [22]), .b(\eq_47_3/LTV [22]), 
        .out(\eq_47_3/LTV2 [22]) );
  nand2 \eq_47_3/ULTI2_22  ( .a(\eq_47_3/LTV1 [22]), .b(\eq_47_3/LTV2 [22]), 
        .out(\eq_47_3/LTV [23]) );
  xor2 \eq_47_3/UEQI_23  ( .a(current_floor_output_elevator2[23]), .b(
        destination_floor_elevator2[23]), .out(n2383) );
  nand2 \eq_47_3/UGTI0_23  ( .a(n2382), .b(current_floor_output_elevator2[23]), 
        .out(\eq_47_3/GTV1 [23]) );
  nand2 \eq_47_3/UGTI1_23  ( .a(\eq_47_3/AEQB [23]), .b(\eq_47_3/GTV [23]), 
        .out(\eq_47_3/GTV2 [23]) );
  nand2 \eq_47_3/UGTI2_23  ( .a(\eq_47_3/GTV1 [23]), .b(\eq_47_3/GTV2 [23]), 
        .out(\eq_47_3/GTV [24]) );
  nand2 \eq_47_3/ULTI0_23  ( .a(n2381), .b(destination_floor_elevator2[23]), 
        .out(\eq_47_3/LTV1 [23]) );
  nand2 \eq_47_3/ULTI1_23  ( .a(\eq_47_3/AEQB [23]), .b(\eq_47_3/LTV [23]), 
        .out(\eq_47_3/LTV2 [23]) );
  nand2 \eq_47_3/ULTI2_23  ( .a(\eq_47_3/LTV1 [23]), .b(\eq_47_3/LTV2 [23]), 
        .out(\eq_47_3/LTV [24]) );
  xor2 \eq_47_3/UEQI_24  ( .a(current_floor_output_elevator2[24]), .b(
        destination_floor_elevator2[24]), .out(n2380) );
  nand2 \eq_47_3/UGTI0_24  ( .a(n2379), .b(current_floor_output_elevator2[24]), 
        .out(\eq_47_3/GTV1 [24]) );
  nand2 \eq_47_3/UGTI1_24  ( .a(\eq_47_3/AEQB [24]), .b(\eq_47_3/GTV [24]), 
        .out(\eq_47_3/GTV2 [24]) );
  nand2 \eq_47_3/UGTI2_24  ( .a(\eq_47_3/GTV1 [24]), .b(\eq_47_3/GTV2 [24]), 
        .out(\eq_47_3/GTV [25]) );
  nand2 \eq_47_3/ULTI0_24  ( .a(n2378), .b(destination_floor_elevator2[24]), 
        .out(\eq_47_3/LTV1 [24]) );
  nand2 \eq_47_3/ULTI1_24  ( .a(\eq_47_3/AEQB [24]), .b(\eq_47_3/LTV [24]), 
        .out(\eq_47_3/LTV2 [24]) );
  nand2 \eq_47_3/ULTI2_24  ( .a(\eq_47_3/LTV1 [24]), .b(\eq_47_3/LTV2 [24]), 
        .out(\eq_47_3/LTV [25]) );
  xor2 \eq_47_3/UEQI_25  ( .a(current_floor_output_elevator2[25]), .b(
        destination_floor_elevator2[25]), .out(n2377) );
  nand2 \eq_47_3/UGTI0_25  ( .a(n2376), .b(current_floor_output_elevator2[25]), 
        .out(\eq_47_3/GTV1 [25]) );
  nand2 \eq_47_3/UGTI1_25  ( .a(\eq_47_3/AEQB [25]), .b(\eq_47_3/GTV [25]), 
        .out(\eq_47_3/GTV2 [25]) );
  nand2 \eq_47_3/UGTI2_25  ( .a(\eq_47_3/GTV1 [25]), .b(\eq_47_3/GTV2 [25]), 
        .out(\eq_47_3/GTV [26]) );
  nand2 \eq_47_3/ULTI0_25  ( .a(n2375), .b(destination_floor_elevator2[25]), 
        .out(\eq_47_3/LTV1 [25]) );
  nand2 \eq_47_3/ULTI1_25  ( .a(\eq_47_3/AEQB [25]), .b(\eq_47_3/LTV [25]), 
        .out(\eq_47_3/LTV2 [25]) );
  nand2 \eq_47_3/ULTI2_25  ( .a(\eq_47_3/LTV1 [25]), .b(\eq_47_3/LTV2 [25]), 
        .out(\eq_47_3/LTV [26]) );
  xor2 \eq_47_3/UEQI_26  ( .a(current_floor_output_elevator2[26]), .b(
        destination_floor_elevator2[26]), .out(n2374) );
  nand2 \eq_47_3/UGTI0_26  ( .a(n2373), .b(current_floor_output_elevator2[26]), 
        .out(\eq_47_3/GTV1 [26]) );
  nand2 \eq_47_3/UGTI1_26  ( .a(\eq_47_3/AEQB [26]), .b(\eq_47_3/GTV [26]), 
        .out(\eq_47_3/GTV2 [26]) );
  nand2 \eq_47_3/UGTI2_26  ( .a(\eq_47_3/GTV1 [26]), .b(\eq_47_3/GTV2 [26]), 
        .out(\eq_47_3/GTV [27]) );
  nand2 \eq_47_3/ULTI0_26  ( .a(n2372), .b(destination_floor_elevator2[26]), 
        .out(\eq_47_3/LTV1 [26]) );
  nand2 \eq_47_3/ULTI1_26  ( .a(\eq_47_3/AEQB [26]), .b(\eq_47_3/LTV [26]), 
        .out(\eq_47_3/LTV2 [26]) );
  nand2 \eq_47_3/ULTI2_26  ( .a(\eq_47_3/LTV1 [26]), .b(\eq_47_3/LTV2 [26]), 
        .out(\eq_47_3/LTV [27]) );
  xor2 \eq_47_3/UEQI_27  ( .a(current_floor_output_elevator2[27]), .b(
        destination_floor_elevator2[27]), .out(n2371) );
  nand2 \eq_47_3/UGTI0_27  ( .a(n2370), .b(current_floor_output_elevator2[27]), 
        .out(\eq_47_3/GTV1 [27]) );
  nand2 \eq_47_3/UGTI1_27  ( .a(\eq_47_3/AEQB [27]), .b(\eq_47_3/GTV [27]), 
        .out(\eq_47_3/GTV2 [27]) );
  nand2 \eq_47_3/UGTI2_27  ( .a(\eq_47_3/GTV1 [27]), .b(\eq_47_3/GTV2 [27]), 
        .out(\eq_47_3/GTV [28]) );
  nand2 \eq_47_3/ULTI0_27  ( .a(n2369), .b(destination_floor_elevator2[27]), 
        .out(\eq_47_3/LTV1 [27]) );
  nand2 \eq_47_3/ULTI1_27  ( .a(\eq_47_3/AEQB [27]), .b(\eq_47_3/LTV [27]), 
        .out(\eq_47_3/LTV2 [27]) );
  nand2 \eq_47_3/ULTI2_27  ( .a(\eq_47_3/LTV1 [27]), .b(\eq_47_3/LTV2 [27]), 
        .out(\eq_47_3/LTV [28]) );
  xor2 \eq_47_3/UEQI_28  ( .a(current_floor_output_elevator2[28]), .b(
        destination_floor_elevator2[28]), .out(n2368) );
  nand2 \eq_47_3/UGTI0_28  ( .a(n2367), .b(current_floor_output_elevator2[28]), 
        .out(\eq_47_3/GTV1 [28]) );
  nand2 \eq_47_3/UGTI1_28  ( .a(\eq_47_3/AEQB [28]), .b(\eq_47_3/GTV [28]), 
        .out(\eq_47_3/GTV2 [28]) );
  nand2 \eq_47_3/UGTI2_28  ( .a(\eq_47_3/GTV1 [28]), .b(\eq_47_3/GTV2 [28]), 
        .out(\eq_47_3/GTV [29]) );
  nand2 \eq_47_3/ULTI0_28  ( .a(n2366), .b(destination_floor_elevator2[28]), 
        .out(\eq_47_3/LTV1 [28]) );
  nand2 \eq_47_3/ULTI1_28  ( .a(\eq_47_3/AEQB [28]), .b(\eq_47_3/LTV [28]), 
        .out(\eq_47_3/LTV2 [28]) );
  nand2 \eq_47_3/ULTI2_28  ( .a(\eq_47_3/LTV1 [28]), .b(\eq_47_3/LTV2 [28]), 
        .out(\eq_47_3/LTV [29]) );
  xor2 \eq_47_3/UEQI_29  ( .a(current_floor_output_elevator2[29]), .b(
        destination_floor_elevator2[29]), .out(n2365) );
  nand2 \eq_47_3/UGTI0_29  ( .a(n2364), .b(current_floor_output_elevator2[29]), 
        .out(\eq_47_3/GTV1 [29]) );
  nand2 \eq_47_3/UGTI1_29  ( .a(\eq_47_3/AEQB [29]), .b(\eq_47_3/GTV [29]), 
        .out(\eq_47_3/GTV2 [29]) );
  nand2 \eq_47_3/UGTI2_29  ( .a(\eq_47_3/GTV1 [29]), .b(\eq_47_3/GTV2 [29]), 
        .out(\eq_47_3/GTV [30]) );
  nand2 \eq_47_3/ULTI0_29  ( .a(n2363), .b(destination_floor_elevator2[29]), 
        .out(\eq_47_3/LTV1 [29]) );
  nand2 \eq_47_3/ULTI1_29  ( .a(\eq_47_3/AEQB [29]), .b(\eq_47_3/LTV [29]), 
        .out(\eq_47_3/LTV2 [29]) );
  nand2 \eq_47_3/ULTI2_29  ( .a(\eq_47_3/LTV1 [29]), .b(\eq_47_3/LTV2 [29]), 
        .out(\eq_47_3/LTV [30]) );
  xor2 \eq_47_3/UEQI_30  ( .a(current_floor_output_elevator2[30]), .b(
        destination_floor_elevator2[30]), .out(n2362) );
  nand2 \eq_47_3/UGTI0_30  ( .a(n2361), .b(current_floor_output_elevator2[30]), 
        .out(\eq_47_3/GTV1 [30]) );
  nand2 \eq_47_3/UGTI1_30  ( .a(\eq_47_3/AEQB [30]), .b(\eq_47_3/GTV [30]), 
        .out(\eq_47_3/GTV2 [30]) );
  nand2 \eq_47_3/UGTI2_30  ( .a(\eq_47_3/GTV1 [30]), .b(\eq_47_3/GTV2 [30]), 
        .out(\eq_47_3/GTV [31]) );
  nand2 \eq_47_3/ULTI0_30  ( .a(n2360), .b(destination_floor_elevator2[30]), 
        .out(\eq_47_3/LTV1 [30]) );
  nand2 \eq_47_3/ULTI1_30  ( .a(\eq_47_3/AEQB [30]), .b(\eq_47_3/LTV [30]), 
        .out(\eq_47_3/LTV2 [30]) );
  nand2 \eq_47_3/ULTI2_30  ( .a(\eq_47_3/LTV1 [30]), .b(\eq_47_3/LTV2 [30]), 
        .out(\eq_47_3/LTV [31]) );
  xor2 \eq_47_3/UEQI_31  ( .a(current_floor_output_elevator2[31]), .b(
        destination_floor_elevator2[31]), .out(n2359) );
  nand2 \eq_47_3/UGTI0_31  ( .a(n2358), .b(current_floor_output_elevator2[31]), 
        .out(\eq_47_3/GTV1 [31]) );
  nand2 \eq_47_3/UGTI1_31  ( .a(\eq_47_3/AEQB [31]), .b(\eq_47_3/GTV [31]), 
        .out(\eq_47_3/GTV2 [31]) );
  nand2 \eq_47_3/UGTI2_31  ( .a(\eq_47_3/GTV1 [31]), .b(\eq_47_3/GTV2 [31]), 
        .out(\eq_47_3/GTV [32]) );
  nand2 \eq_47_3/ULTI0_31  ( .a(n2357), .b(destination_floor_elevator2[31]), 
        .out(\eq_47_3/LTV1 [31]) );
  nand2 \eq_47_3/ULTI1_31  ( .a(\eq_47_3/AEQB [31]), .b(\eq_47_3/LTV [31]), 
        .out(\eq_47_3/LTV2 [31]) );
  nand2 \eq_47_3/ULTI2_31  ( .a(\eq_47_3/LTV1 [31]), .b(\eq_47_3/LTV2 [31]), 
        .out(\eq_47_3/LTV [32]) );
  xor2 \eq_47_3/UEQI_32  ( .a(current_floor_output_elevator2[32]), .b(
        destination_floor_elevator2[32]), .out(n2356) );
  nand2 \eq_47_3/UGTI0_32  ( .a(n2355), .b(current_floor_output_elevator2[32]), 
        .out(\eq_47_3/GTV1 [32]) );
  nand2 \eq_47_3/UGTI1_32  ( .a(\eq_47_3/AEQB [32]), .b(\eq_47_3/GTV [32]), 
        .out(\eq_47_3/GTV2 [32]) );
  nand2 \eq_47_3/UGTI2_32  ( .a(\eq_47_3/GTV1 [32]), .b(\eq_47_3/GTV2 [32]), 
        .out(\eq_47_3/GTV [33]) );
  nand2 \eq_47_3/ULTI0_32  ( .a(n2354), .b(destination_floor_elevator2[32]), 
        .out(\eq_47_3/LTV1 [32]) );
  nand2 \eq_47_3/ULTI1_32  ( .a(\eq_47_3/AEQB [32]), .b(\eq_47_3/LTV [32]), 
        .out(\eq_47_3/LTV2 [32]) );
  nand2 \eq_47_3/ULTI2_32  ( .a(\eq_47_3/LTV1 [32]), .b(\eq_47_3/LTV2 [32]), 
        .out(\eq_47_3/LTV [33]) );
  xor2 \eq_47_3/UEQI_33  ( .a(current_floor_output_elevator2[33]), .b(
        destination_floor_elevator2[33]), .out(n2353) );
  nand2 \eq_47_3/UGTI0_33  ( .a(n2352), .b(current_floor_output_elevator2[33]), 
        .out(\eq_47_3/GTV1 [33]) );
  nand2 \eq_47_3/UGTI1_33  ( .a(\eq_47_3/AEQB [33]), .b(\eq_47_3/GTV [33]), 
        .out(\eq_47_3/GTV2 [33]) );
  nand2 \eq_47_3/UGTI2_33  ( .a(\eq_47_3/GTV1 [33]), .b(\eq_47_3/GTV2 [33]), 
        .out(\eq_47_3/GTV [34]) );
  nand2 \eq_47_3/ULTI0_33  ( .a(n2351), .b(destination_floor_elevator2[33]), 
        .out(\eq_47_3/LTV1 [33]) );
  nand2 \eq_47_3/ULTI1_33  ( .a(\eq_47_3/AEQB [33]), .b(\eq_47_3/LTV [33]), 
        .out(\eq_47_3/LTV2 [33]) );
  nand2 \eq_47_3/ULTI2_33  ( .a(\eq_47_3/LTV1 [33]), .b(\eq_47_3/LTV2 [33]), 
        .out(\eq_47_3/LTV [34]) );
  xor2 \eq_47_3/UEQI_34  ( .a(current_floor_output_elevator2[34]), .b(
        destination_floor_elevator2[34]), .out(n2350) );
  nand2 \eq_47_3/UGTI0_34  ( .a(n2349), .b(current_floor_output_elevator2[34]), 
        .out(\eq_47_3/GTV1 [34]) );
  nand2 \eq_47_3/UGTI1_34  ( .a(\eq_47_3/AEQB [34]), .b(\eq_47_3/GTV [34]), 
        .out(\eq_47_3/GTV2 [34]) );
  nand2 \eq_47_3/UGTI2_34  ( .a(\eq_47_3/GTV1 [34]), .b(\eq_47_3/GTV2 [34]), 
        .out(\eq_47_3/GTV [35]) );
  nand2 \eq_47_3/ULTI0_34  ( .a(n2348), .b(destination_floor_elevator2[34]), 
        .out(\eq_47_3/LTV1 [34]) );
  nand2 \eq_47_3/ULTI1_34  ( .a(\eq_47_3/AEQB [34]), .b(\eq_47_3/LTV [34]), 
        .out(\eq_47_3/LTV2 [34]) );
  nand2 \eq_47_3/ULTI2_34  ( .a(\eq_47_3/LTV1 [34]), .b(\eq_47_3/LTV2 [34]), 
        .out(\eq_47_3/LTV [35]) );
  xor2 \eq_47_3/UEQI_35  ( .a(current_floor_output_elevator2[35]), .b(
        destination_floor_elevator2[35]), .out(n2347) );
  nand2 \eq_47_3/UGTI0_35  ( .a(n2346), .b(current_floor_output_elevator2[35]), 
        .out(\eq_47_3/GTV1 [35]) );
  nand2 \eq_47_3/UGTI1_35  ( .a(\eq_47_3/AEQB [35]), .b(\eq_47_3/GTV [35]), 
        .out(\eq_47_3/GTV2 [35]) );
  nand2 \eq_47_3/UGTI2_35  ( .a(\eq_47_3/GTV1 [35]), .b(\eq_47_3/GTV2 [35]), 
        .out(\eq_47_3/GTV [36]) );
  nand2 \eq_47_3/ULTI0_35  ( .a(n2345), .b(destination_floor_elevator2[35]), 
        .out(\eq_47_3/LTV1 [35]) );
  nand2 \eq_47_3/ULTI1_35  ( .a(\eq_47_3/AEQB [35]), .b(\eq_47_3/LTV [35]), 
        .out(\eq_47_3/LTV2 [35]) );
  nand2 \eq_47_3/ULTI2_35  ( .a(\eq_47_3/LTV1 [35]), .b(\eq_47_3/LTV2 [35]), 
        .out(\eq_47_3/LTV [36]) );
  xor2 \eq_47_3/UEQI_36  ( .a(current_floor_output_elevator2[36]), .b(
        destination_floor_elevator2[36]), .out(n2344) );
  nand2 \eq_47_3/UGTI0_36  ( .a(n2343), .b(current_floor_output_elevator2[36]), 
        .out(\eq_47_3/GTV1 [36]) );
  nand2 \eq_47_3/UGTI1_36  ( .a(\eq_47_3/AEQB [36]), .b(\eq_47_3/GTV [36]), 
        .out(\eq_47_3/GTV2 [36]) );
  nand2 \eq_47_3/UGTI2_36  ( .a(\eq_47_3/GTV1 [36]), .b(\eq_47_3/GTV2 [36]), 
        .out(\eq_47_3/GTV [37]) );
  nand2 \eq_47_3/ULTI0_36  ( .a(n2342), .b(destination_floor_elevator2[36]), 
        .out(\eq_47_3/LTV1 [36]) );
  nand2 \eq_47_3/ULTI1_36  ( .a(\eq_47_3/AEQB [36]), .b(\eq_47_3/LTV [36]), 
        .out(\eq_47_3/LTV2 [36]) );
  nand2 \eq_47_3/ULTI2_36  ( .a(\eq_47_3/LTV1 [36]), .b(\eq_47_3/LTV2 [36]), 
        .out(\eq_47_3/LTV [37]) );
  xor2 \eq_47_3/UEQI_37  ( .a(current_floor_output_elevator2[37]), .b(
        destination_floor_elevator2[37]), .out(n2341) );
  nand2 \eq_47_3/UGTI0_37  ( .a(n2340), .b(current_floor_output_elevator2[37]), 
        .out(\eq_47_3/GTV1 [37]) );
  nand2 \eq_47_3/UGTI1_37  ( .a(\eq_47_3/AEQB [37]), .b(\eq_47_3/GTV [37]), 
        .out(\eq_47_3/GTV2 [37]) );
  nand2 \eq_47_3/UGTI2_37  ( .a(\eq_47_3/GTV1 [37]), .b(\eq_47_3/GTV2 [37]), 
        .out(\eq_47_3/GTV [38]) );
  nand2 \eq_47_3/ULTI0_37  ( .a(n2339), .b(destination_floor_elevator2[37]), 
        .out(\eq_47_3/LTV1 [37]) );
  nand2 \eq_47_3/ULTI1_37  ( .a(\eq_47_3/AEQB [37]), .b(\eq_47_3/LTV [37]), 
        .out(\eq_47_3/LTV2 [37]) );
  nand2 \eq_47_3/ULTI2_37  ( .a(\eq_47_3/LTV1 [37]), .b(\eq_47_3/LTV2 [37]), 
        .out(\eq_47_3/LTV [38]) );
  xor2 \eq_47_3/UEQI_38  ( .a(current_floor_output_elevator2[38]), .b(
        destination_floor_elevator2[38]), .out(n2338) );
  nand2 \eq_47_3/UGTI0_38  ( .a(n2337), .b(current_floor_output_elevator2[38]), 
        .out(\eq_47_3/GTV1 [38]) );
  nand2 \eq_47_3/UGTI1_38  ( .a(\eq_47_3/AEQB [38]), .b(\eq_47_3/GTV [38]), 
        .out(\eq_47_3/GTV2 [38]) );
  nand2 \eq_47_3/UGTI2_38  ( .a(\eq_47_3/GTV1 [38]), .b(\eq_47_3/GTV2 [38]), 
        .out(\eq_47_3/GTV [39]) );
  nand2 \eq_47_3/ULTI0_38  ( .a(n2336), .b(destination_floor_elevator2[38]), 
        .out(\eq_47_3/LTV1 [38]) );
  nand2 \eq_47_3/ULTI1_38  ( .a(\eq_47_3/AEQB [38]), .b(\eq_47_3/LTV [38]), 
        .out(\eq_47_3/LTV2 [38]) );
  nand2 \eq_47_3/ULTI2_38  ( .a(\eq_47_3/LTV1 [38]), .b(\eq_47_3/LTV2 [38]), 
        .out(\eq_47_3/LTV [39]) );
  xor2 \eq_47_3/UEQI_39  ( .a(current_floor_output_elevator2[39]), .b(
        destination_floor_elevator2[39]), .out(n2335) );
  nand2 \eq_47_3/UGTI0_39  ( .a(n2334), .b(current_floor_output_elevator2[39]), 
        .out(\eq_47_3/GTV1 [39]) );
  nand2 \eq_47_3/UGTI1_39  ( .a(\eq_47_3/AEQB [39]), .b(\eq_47_3/GTV [39]), 
        .out(\eq_47_3/GTV2 [39]) );
  nand2 \eq_47_3/UGTI2_39  ( .a(\eq_47_3/GTV1 [39]), .b(\eq_47_3/GTV2 [39]), 
        .out(\eq_47_3/GTV [40]) );
  nand2 \eq_47_3/ULTI0_39  ( .a(n2333), .b(destination_floor_elevator2[39]), 
        .out(\eq_47_3/LTV1 [39]) );
  nand2 \eq_47_3/ULTI1_39  ( .a(\eq_47_3/AEQB [39]), .b(\eq_47_3/LTV [39]), 
        .out(\eq_47_3/LTV2 [39]) );
  nand2 \eq_47_3/ULTI2_39  ( .a(\eq_47_3/LTV1 [39]), .b(\eq_47_3/LTV2 [39]), 
        .out(\eq_47_3/LTV [40]) );
  xor2 \eq_47_3/UEQI_40  ( .a(current_floor_output_elevator2[40]), .b(
        destination_floor_elevator2[40]), .out(n2332) );
  nand2 \eq_47_3/UGTI0_40  ( .a(n2331), .b(current_floor_output_elevator2[40]), 
        .out(\eq_47_3/GTV1 [40]) );
  nand2 \eq_47_3/UGTI1_40  ( .a(\eq_47_3/AEQB [40]), .b(\eq_47_3/GTV [40]), 
        .out(\eq_47_3/GTV2 [40]) );
  nand2 \eq_47_3/UGTI2_40  ( .a(\eq_47_3/GTV1 [40]), .b(\eq_47_3/GTV2 [40]), 
        .out(\eq_47_3/GTV [41]) );
  nand2 \eq_47_3/ULTI0_40  ( .a(n2330), .b(destination_floor_elevator2[40]), 
        .out(\eq_47_3/LTV1 [40]) );
  nand2 \eq_47_3/ULTI1_40  ( .a(\eq_47_3/AEQB [40]), .b(\eq_47_3/LTV [40]), 
        .out(\eq_47_3/LTV2 [40]) );
  nand2 \eq_47_3/ULTI2_40  ( .a(\eq_47_3/LTV1 [40]), .b(\eq_47_3/LTV2 [40]), 
        .out(\eq_47_3/LTV [41]) );
  xor2 \eq_47_3/UEQI_41  ( .a(current_floor_output_elevator2[41]), .b(
        destination_floor_elevator2[41]), .out(n2329) );
  nand2 \eq_47_3/UGTI0_41  ( .a(n2328), .b(current_floor_output_elevator2[41]), 
        .out(\eq_47_3/GTV1 [41]) );
  nand2 \eq_47_3/UGTI1_41  ( .a(\eq_47_3/AEQB [41]), .b(\eq_47_3/GTV [41]), 
        .out(\eq_47_3/GTV2 [41]) );
  nand2 \eq_47_3/UGTI2_41  ( .a(\eq_47_3/GTV1 [41]), .b(\eq_47_3/GTV2 [41]), 
        .out(\eq_47_3/GTV [42]) );
  nand2 \eq_47_3/ULTI0_41  ( .a(n2327), .b(destination_floor_elevator2[41]), 
        .out(\eq_47_3/LTV1 [41]) );
  nand2 \eq_47_3/ULTI1_41  ( .a(\eq_47_3/AEQB [41]), .b(\eq_47_3/LTV [41]), 
        .out(\eq_47_3/LTV2 [41]) );
  nand2 \eq_47_3/ULTI2_41  ( .a(\eq_47_3/LTV1 [41]), .b(\eq_47_3/LTV2 [41]), 
        .out(\eq_47_3/LTV [42]) );
  xor2 \eq_47_3/UEQI_42  ( .a(current_floor_output_elevator2[42]), .b(
        destination_floor_elevator2[42]), .out(n2326) );
  nand2 \eq_47_3/UGTI0_42  ( .a(n2325), .b(current_floor_output_elevator2[42]), 
        .out(\eq_47_3/GTV1 [42]) );
  nand2 \eq_47_3/UGTI1_42  ( .a(\eq_47_3/AEQB [42]), .b(\eq_47_3/GTV [42]), 
        .out(\eq_47_3/GTV2 [42]) );
  nand2 \eq_47_3/UGTI2_42  ( .a(\eq_47_3/GTV1 [42]), .b(\eq_47_3/GTV2 [42]), 
        .out(\eq_47_3/GTV [43]) );
  nand2 \eq_47_3/ULTI0_42  ( .a(n2324), .b(destination_floor_elevator2[42]), 
        .out(\eq_47_3/LTV1 [42]) );
  nand2 \eq_47_3/ULTI1_42  ( .a(\eq_47_3/AEQB [42]), .b(\eq_47_3/LTV [42]), 
        .out(\eq_47_3/LTV2 [42]) );
  nand2 \eq_47_3/ULTI2_42  ( .a(\eq_47_3/LTV1 [42]), .b(\eq_47_3/LTV2 [42]), 
        .out(\eq_47_3/LTV [43]) );
  xor2 \eq_47_3/UEQI_43  ( .a(current_floor_output_elevator2[43]), .b(
        destination_floor_elevator2[43]), .out(n2323) );
  nand2 \eq_47_3/UGTI0_43  ( .a(n2322), .b(current_floor_output_elevator2[43]), 
        .out(\eq_47_3/GTV1 [43]) );
  nand2 \eq_47_3/UGTI1_43  ( .a(\eq_47_3/AEQB [43]), .b(\eq_47_3/GTV [43]), 
        .out(\eq_47_3/GTV2 [43]) );
  nand2 \eq_47_3/UGTI2_43  ( .a(\eq_47_3/GTV1 [43]), .b(\eq_47_3/GTV2 [43]), 
        .out(\eq_47_3/GTV [44]) );
  nand2 \eq_47_3/ULTI0_43  ( .a(n2321), .b(destination_floor_elevator2[43]), 
        .out(\eq_47_3/LTV1 [43]) );
  nand2 \eq_47_3/ULTI1_43  ( .a(\eq_47_3/AEQB [43]), .b(\eq_47_3/LTV [43]), 
        .out(\eq_47_3/LTV2 [43]) );
  nand2 \eq_47_3/ULTI2_43  ( .a(\eq_47_3/LTV1 [43]), .b(\eq_47_3/LTV2 [43]), 
        .out(\eq_47_3/LTV [44]) );
  xor2 \eq_47_3/UEQI_44  ( .a(current_floor_output_elevator2[44]), .b(
        destination_floor_elevator2[44]), .out(n2320) );
  nand2 \eq_47_3/UGTI0_44  ( .a(n2319), .b(current_floor_output_elevator2[44]), 
        .out(\eq_47_3/GTV1 [44]) );
  nand2 \eq_47_3/UGTI1_44  ( .a(\eq_47_3/AEQB [44]), .b(\eq_47_3/GTV [44]), 
        .out(\eq_47_3/GTV2 [44]) );
  nand2 \eq_47_3/UGTI2_44  ( .a(\eq_47_3/GTV1 [44]), .b(\eq_47_3/GTV2 [44]), 
        .out(\eq_47_3/GTV [45]) );
  nand2 \eq_47_3/ULTI0_44  ( .a(n2318), .b(destination_floor_elevator2[44]), 
        .out(\eq_47_3/LTV1 [44]) );
  nand2 \eq_47_3/ULTI1_44  ( .a(\eq_47_3/AEQB [44]), .b(\eq_47_3/LTV [44]), 
        .out(\eq_47_3/LTV2 [44]) );
  nand2 \eq_47_3/ULTI2_44  ( .a(\eq_47_3/LTV1 [44]), .b(\eq_47_3/LTV2 [44]), 
        .out(\eq_47_3/LTV [45]) );
  xor2 \eq_47_3/UEQI_45  ( .a(current_floor_output_elevator2[45]), .b(
        destination_floor_elevator2[45]), .out(n2317) );
  nand2 \eq_47_3/UGTI0_45  ( .a(n2316), .b(current_floor_output_elevator2[45]), 
        .out(\eq_47_3/GTV1 [45]) );
  nand2 \eq_47_3/UGTI1_45  ( .a(\eq_47_3/AEQB [45]), .b(\eq_47_3/GTV [45]), 
        .out(\eq_47_3/GTV2 [45]) );
  nand2 \eq_47_3/UGTI2_45  ( .a(\eq_47_3/GTV1 [45]), .b(\eq_47_3/GTV2 [45]), 
        .out(\eq_47_3/GTV [46]) );
  nand2 \eq_47_3/ULTI0_45  ( .a(n2315), .b(destination_floor_elevator2[45]), 
        .out(\eq_47_3/LTV1 [45]) );
  nand2 \eq_47_3/ULTI1_45  ( .a(\eq_47_3/AEQB [45]), .b(\eq_47_3/LTV [45]), 
        .out(\eq_47_3/LTV2 [45]) );
  nand2 \eq_47_3/ULTI2_45  ( .a(\eq_47_3/LTV1 [45]), .b(\eq_47_3/LTV2 [45]), 
        .out(\eq_47_3/LTV [46]) );
  xor2 \eq_47_3/UEQI_46  ( .a(current_floor_output_elevator2[46]), .b(
        destination_floor_elevator2[46]), .out(n2314) );
  nand2 \eq_47_3/UGTI0_46  ( .a(n2313), .b(current_floor_output_elevator2[46]), 
        .out(\eq_47_3/GTV1 [46]) );
  nand2 \eq_47_3/UGTI1_46  ( .a(\eq_47_3/AEQB [46]), .b(\eq_47_3/GTV [46]), 
        .out(\eq_47_3/GTV2 [46]) );
  nand2 \eq_47_3/UGTI2_46  ( .a(\eq_47_3/GTV1 [46]), .b(\eq_47_3/GTV2 [46]), 
        .out(\eq_47_3/GTV [47]) );
  nand2 \eq_47_3/ULTI0_46  ( .a(n2312), .b(destination_floor_elevator2[46]), 
        .out(\eq_47_3/LTV1 [46]) );
  nand2 \eq_47_3/ULTI1_46  ( .a(\eq_47_3/AEQB [46]), .b(\eq_47_3/LTV [46]), 
        .out(\eq_47_3/LTV2 [46]) );
  nand2 \eq_47_3/ULTI2_46  ( .a(\eq_47_3/LTV1 [46]), .b(\eq_47_3/LTV2 [46]), 
        .out(\eq_47_3/LTV [47]) );
  xor2 \eq_47_3/UEQI_47  ( .a(current_floor_output_elevator2[47]), .b(
        destination_floor_elevator2[47]), .out(n2311) );
  nand2 \eq_47_3/UGTI0_47  ( .a(n2310), .b(current_floor_output_elevator2[47]), 
        .out(\eq_47_3/GTV1 [47]) );
  nand2 \eq_47_3/UGTI1_47  ( .a(\eq_47_3/AEQB [47]), .b(\eq_47_3/GTV [47]), 
        .out(\eq_47_3/GTV2 [47]) );
  nand2 \eq_47_3/UGTI2_47  ( .a(\eq_47_3/GTV1 [47]), .b(\eq_47_3/GTV2 [47]), 
        .out(\eq_47_3/GTV [48]) );
  nand2 \eq_47_3/ULTI0_47  ( .a(n2309), .b(destination_floor_elevator2[47]), 
        .out(\eq_47_3/LTV1 [47]) );
  nand2 \eq_47_3/ULTI1_47  ( .a(\eq_47_3/AEQB [47]), .b(\eq_47_3/LTV [47]), 
        .out(\eq_47_3/LTV2 [47]) );
  nand2 \eq_47_3/ULTI2_47  ( .a(\eq_47_3/LTV1 [47]), .b(\eq_47_3/LTV2 [47]), 
        .out(\eq_47_3/LTV [48]) );
  xor2 \eq_47_3/UEQI_48  ( .a(current_floor_output_elevator2[48]), .b(
        destination_floor_elevator2[48]), .out(n2308) );
  nand2 \eq_47_3/UGTI0_48  ( .a(n2307), .b(current_floor_output_elevator2[48]), 
        .out(\eq_47_3/GTV1 [48]) );
  nand2 \eq_47_3/UGTI1_48  ( .a(\eq_47_3/AEQB [48]), .b(\eq_47_3/GTV [48]), 
        .out(\eq_47_3/GTV2 [48]) );
  nand2 \eq_47_3/UGTI2_48  ( .a(\eq_47_3/GTV1 [48]), .b(\eq_47_3/GTV2 [48]), 
        .out(\eq_47_3/GTV [49]) );
  nand2 \eq_47_3/ULTI0_48  ( .a(n2306), .b(destination_floor_elevator2[48]), 
        .out(\eq_47_3/LTV1 [48]) );
  nand2 \eq_47_3/ULTI1_48  ( .a(\eq_47_3/AEQB [48]), .b(\eq_47_3/LTV [48]), 
        .out(\eq_47_3/LTV2 [48]) );
  nand2 \eq_47_3/ULTI2_48  ( .a(\eq_47_3/LTV1 [48]), .b(\eq_47_3/LTV2 [48]), 
        .out(\eq_47_3/LTV [49]) );
  xor2 \eq_47_3/UEQI_49  ( .a(current_floor_output_elevator2[49]), .b(
        destination_floor_elevator2[49]), .out(n2305) );
  nand2 \eq_47_3/UGTI0_49  ( .a(n2304), .b(current_floor_output_elevator2[49]), 
        .out(\eq_47_3/GTV1 [49]) );
  nand2 \eq_47_3/UGTI1_49  ( .a(\eq_47_3/AEQB [49]), .b(\eq_47_3/GTV [49]), 
        .out(\eq_47_3/GTV2 [49]) );
  nand2 \eq_47_3/UGTI2_49  ( .a(\eq_47_3/GTV1 [49]), .b(\eq_47_3/GTV2 [49]), 
        .out(\eq_47_3/GTV [50]) );
  nand2 \eq_47_3/ULTI0_49  ( .a(n2303), .b(destination_floor_elevator2[49]), 
        .out(\eq_47_3/LTV1 [49]) );
  nand2 \eq_47_3/ULTI1_49  ( .a(\eq_47_3/AEQB [49]), .b(\eq_47_3/LTV [49]), 
        .out(\eq_47_3/LTV2 [49]) );
  nand2 \eq_47_3/ULTI2_49  ( .a(\eq_47_3/LTV1 [49]), .b(\eq_47_3/LTV2 [49]), 
        .out(\eq_47_3/LTV [50]) );
  xor2 \eq_47_3/UEQI_50  ( .a(current_floor_output_elevator2[50]), .b(
        destination_floor_elevator2[50]), .out(n2302) );
  nand2 \eq_47_3/UGTI0_50  ( .a(n2301), .b(current_floor_output_elevator2[50]), 
        .out(\eq_47_3/GTV1 [50]) );
  nand2 \eq_47_3/UGTI1_50  ( .a(\eq_47_3/AEQB [50]), .b(\eq_47_3/GTV [50]), 
        .out(\eq_47_3/GTV2 [50]) );
  nand2 \eq_47_3/UGTI2_50  ( .a(\eq_47_3/GTV1 [50]), .b(\eq_47_3/GTV2 [50]), 
        .out(\eq_47_3/GTV [51]) );
  nand2 \eq_47_3/ULTI0_50  ( .a(n2300), .b(destination_floor_elevator2[50]), 
        .out(\eq_47_3/LTV1 [50]) );
  nand2 \eq_47_3/ULTI1_50  ( .a(\eq_47_3/AEQB [50]), .b(\eq_47_3/LTV [50]), 
        .out(\eq_47_3/LTV2 [50]) );
  nand2 \eq_47_3/ULTI2_50  ( .a(\eq_47_3/LTV1 [50]), .b(\eq_47_3/LTV2 [50]), 
        .out(\eq_47_3/LTV [51]) );
  xor2 \eq_47_3/UEQI_51  ( .a(current_floor_output_elevator2[51]), .b(
        destination_floor_elevator2[51]), .out(n2299) );
  nand2 \eq_47_3/UGTI0_51  ( .a(n2298), .b(current_floor_output_elevator2[51]), 
        .out(\eq_47_3/GTV1 [51]) );
  nand2 \eq_47_3/UGTI1_51  ( .a(\eq_47_3/AEQB [51]), .b(\eq_47_3/GTV [51]), 
        .out(\eq_47_3/GTV2 [51]) );
  nand2 \eq_47_3/UGTI2_51  ( .a(\eq_47_3/GTV1 [51]), .b(\eq_47_3/GTV2 [51]), 
        .out(\eq_47_3/GTV [52]) );
  nand2 \eq_47_3/ULTI0_51  ( .a(n2297), .b(destination_floor_elevator2[51]), 
        .out(\eq_47_3/LTV1 [51]) );
  nand2 \eq_47_3/ULTI1_51  ( .a(\eq_47_3/AEQB [51]), .b(\eq_47_3/LTV [51]), 
        .out(\eq_47_3/LTV2 [51]) );
  nand2 \eq_47_3/ULTI2_51  ( .a(\eq_47_3/LTV1 [51]), .b(\eq_47_3/LTV2 [51]), 
        .out(\eq_47_3/LTV [52]) );
  xor2 \eq_47_3/UEQI_52  ( .a(current_floor_output_elevator2[52]), .b(
        destination_floor_elevator2[52]), .out(n2296) );
  nand2 \eq_47_3/UGTI0_52  ( .a(n2295), .b(current_floor_output_elevator2[52]), 
        .out(\eq_47_3/GTV1 [52]) );
  nand2 \eq_47_3/UGTI1_52  ( .a(\eq_47_3/AEQB [52]), .b(\eq_47_3/GTV [52]), 
        .out(\eq_47_3/GTV2 [52]) );
  nand2 \eq_47_3/UGTI2_52  ( .a(\eq_47_3/GTV1 [52]), .b(\eq_47_3/GTV2 [52]), 
        .out(\eq_47_3/GTV [53]) );
  nand2 \eq_47_3/ULTI0_52  ( .a(n2294), .b(destination_floor_elevator2[52]), 
        .out(\eq_47_3/LTV1 [52]) );
  nand2 \eq_47_3/ULTI1_52  ( .a(\eq_47_3/AEQB [52]), .b(\eq_47_3/LTV [52]), 
        .out(\eq_47_3/LTV2 [52]) );
  nand2 \eq_47_3/ULTI2_52  ( .a(\eq_47_3/LTV1 [52]), .b(\eq_47_3/LTV2 [52]), 
        .out(\eq_47_3/LTV [53]) );
  xor2 \eq_47_3/UEQI_53  ( .a(current_floor_output_elevator2[53]), .b(
        destination_floor_elevator2[53]), .out(n2293) );
  nand2 \eq_47_3/UGTI0_53  ( .a(n2292), .b(current_floor_output_elevator2[53]), 
        .out(\eq_47_3/GTV1 [53]) );
  nand2 \eq_47_3/UGTI1_53  ( .a(\eq_47_3/AEQB [53]), .b(\eq_47_3/GTV [53]), 
        .out(\eq_47_3/GTV2 [53]) );
  nand2 \eq_47_3/UGTI2_53  ( .a(\eq_47_3/GTV1 [53]), .b(\eq_47_3/GTV2 [53]), 
        .out(\eq_47_3/GTV [54]) );
  nand2 \eq_47_3/ULTI0_53  ( .a(n2291), .b(destination_floor_elevator2[53]), 
        .out(\eq_47_3/LTV1 [53]) );
  nand2 \eq_47_3/ULTI1_53  ( .a(\eq_47_3/AEQB [53]), .b(\eq_47_3/LTV [53]), 
        .out(\eq_47_3/LTV2 [53]) );
  nand2 \eq_47_3/ULTI2_53  ( .a(\eq_47_3/LTV1 [53]), .b(\eq_47_3/LTV2 [53]), 
        .out(\eq_47_3/LTV [54]) );
  xor2 \eq_47_3/UEQI_54  ( .a(current_floor_output_elevator2[54]), .b(
        destination_floor_elevator2[54]), .out(n2290) );
  nand2 \eq_47_3/UGTI0_54  ( .a(n2289), .b(current_floor_output_elevator2[54]), 
        .out(\eq_47_3/GTV1 [54]) );
  nand2 \eq_47_3/UGTI1_54  ( .a(\eq_47_3/AEQB [54]), .b(\eq_47_3/GTV [54]), 
        .out(\eq_47_3/GTV2 [54]) );
  nand2 \eq_47_3/UGTI2_54  ( .a(\eq_47_3/GTV1 [54]), .b(\eq_47_3/GTV2 [54]), 
        .out(\eq_47_3/GTV [55]) );
  nand2 \eq_47_3/ULTI0_54  ( .a(n2288), .b(destination_floor_elevator2[54]), 
        .out(\eq_47_3/LTV1 [54]) );
  nand2 \eq_47_3/ULTI1_54  ( .a(\eq_47_3/AEQB [54]), .b(\eq_47_3/LTV [54]), 
        .out(\eq_47_3/LTV2 [54]) );
  nand2 \eq_47_3/ULTI2_54  ( .a(\eq_47_3/LTV1 [54]), .b(\eq_47_3/LTV2 [54]), 
        .out(\eq_47_3/LTV [55]) );
  xor2 \eq_47_3/UEQI_55  ( .a(current_floor_output_elevator2[55]), .b(
        destination_floor_elevator2[55]), .out(n2287) );
  nand2 \eq_47_3/UGTI0_55  ( .a(n2286), .b(current_floor_output_elevator2[55]), 
        .out(\eq_47_3/GTV1 [55]) );
  nand2 \eq_47_3/UGTI1_55  ( .a(\eq_47_3/AEQB [55]), .b(\eq_47_3/GTV [55]), 
        .out(\eq_47_3/GTV2 [55]) );
  nand2 \eq_47_3/UGTI2_55  ( .a(\eq_47_3/GTV1 [55]), .b(\eq_47_3/GTV2 [55]), 
        .out(\eq_47_3/GTV [56]) );
  nand2 \eq_47_3/ULTI0_55  ( .a(n2285), .b(destination_floor_elevator2[55]), 
        .out(\eq_47_3/LTV1 [55]) );
  nand2 \eq_47_3/ULTI1_55  ( .a(\eq_47_3/AEQB [55]), .b(\eq_47_3/LTV [55]), 
        .out(\eq_47_3/LTV2 [55]) );
  nand2 \eq_47_3/ULTI2_55  ( .a(\eq_47_3/LTV1 [55]), .b(\eq_47_3/LTV2 [55]), 
        .out(\eq_47_3/LTV [56]) );
  xor2 \eq_47_3/UEQI_56  ( .a(current_floor_output_elevator2[56]), .b(
        destination_floor_elevator2[56]), .out(n2284) );
  nand2 \eq_47_3/UGTI0_56  ( .a(n2283), .b(current_floor_output_elevator2[56]), 
        .out(\eq_47_3/GTV1 [56]) );
  nand2 \eq_47_3/UGTI1_56  ( .a(\eq_47_3/AEQB [56]), .b(\eq_47_3/GTV [56]), 
        .out(\eq_47_3/GTV2 [56]) );
  nand2 \eq_47_3/UGTI2_56  ( .a(\eq_47_3/GTV1 [56]), .b(\eq_47_3/GTV2 [56]), 
        .out(\eq_47_3/GTV [57]) );
  nand2 \eq_47_3/ULTI0_56  ( .a(n2282), .b(destination_floor_elevator2[56]), 
        .out(\eq_47_3/LTV1 [56]) );
  nand2 \eq_47_3/ULTI1_56  ( .a(\eq_47_3/AEQB [56]), .b(\eq_47_3/LTV [56]), 
        .out(\eq_47_3/LTV2 [56]) );
  nand2 \eq_47_3/ULTI2_56  ( .a(\eq_47_3/LTV1 [56]), .b(\eq_47_3/LTV2 [56]), 
        .out(\eq_47_3/LTV [57]) );
  xor2 \eq_47_3/UEQI_57  ( .a(current_floor_output_elevator2[57]), .b(
        destination_floor_elevator2[57]), .out(n2281) );
  nand2 \eq_47_3/UGTI0_57  ( .a(n2280), .b(current_floor_output_elevator2[57]), 
        .out(\eq_47_3/GTV1 [57]) );
  nand2 \eq_47_3/UGTI1_57  ( .a(\eq_47_3/AEQB [57]), .b(\eq_47_3/GTV [57]), 
        .out(\eq_47_3/GTV2 [57]) );
  nand2 \eq_47_3/UGTI2_57  ( .a(\eq_47_3/GTV1 [57]), .b(\eq_47_3/GTV2 [57]), 
        .out(\eq_47_3/GTV [58]) );
  nand2 \eq_47_3/ULTI0_57  ( .a(n2279), .b(destination_floor_elevator2[57]), 
        .out(\eq_47_3/LTV1 [57]) );
  nand2 \eq_47_3/ULTI1_57  ( .a(\eq_47_3/AEQB [57]), .b(\eq_47_3/LTV [57]), 
        .out(\eq_47_3/LTV2 [57]) );
  nand2 \eq_47_3/ULTI2_57  ( .a(\eq_47_3/LTV1 [57]), .b(\eq_47_3/LTV2 [57]), 
        .out(\eq_47_3/LTV [58]) );
  xor2 \eq_47_3/UEQI_58  ( .a(current_floor_output_elevator2[58]), .b(
        destination_floor_elevator2[58]), .out(n2278) );
  nand2 \eq_47_3/UGTI0_58  ( .a(n2277), .b(current_floor_output_elevator2[58]), 
        .out(\eq_47_3/GTV1 [58]) );
  nand2 \eq_47_3/UGTI1_58  ( .a(\eq_47_3/AEQB [58]), .b(\eq_47_3/GTV [58]), 
        .out(\eq_47_3/GTV2 [58]) );
  nand2 \eq_47_3/UGTI2_58  ( .a(\eq_47_3/GTV1 [58]), .b(\eq_47_3/GTV2 [58]), 
        .out(\eq_47_3/GTV [59]) );
  nand2 \eq_47_3/ULTI0_58  ( .a(n2276), .b(destination_floor_elevator2[58]), 
        .out(\eq_47_3/LTV1 [58]) );
  nand2 \eq_47_3/ULTI1_58  ( .a(\eq_47_3/AEQB [58]), .b(\eq_47_3/LTV [58]), 
        .out(\eq_47_3/LTV2 [58]) );
  nand2 \eq_47_3/ULTI2_58  ( .a(\eq_47_3/LTV1 [58]), .b(\eq_47_3/LTV2 [58]), 
        .out(\eq_47_3/LTV [59]) );
  xor2 \eq_47_3/UEQI_59  ( .a(current_floor_output_elevator2[59]), .b(
        destination_floor_elevator2[59]), .out(n2275) );
  nand2 \eq_47_3/UGTI0_59  ( .a(n2274), .b(current_floor_output_elevator2[59]), 
        .out(\eq_47_3/GTV1 [59]) );
  nand2 \eq_47_3/UGTI1_59  ( .a(\eq_47_3/AEQB [59]), .b(\eq_47_3/GTV [59]), 
        .out(\eq_47_3/GTV2 [59]) );
  nand2 \eq_47_3/UGTI2_59  ( .a(\eq_47_3/GTV1 [59]), .b(\eq_47_3/GTV2 [59]), 
        .out(\eq_47_3/GTV [60]) );
  nand2 \eq_47_3/ULTI0_59  ( .a(n2273), .b(destination_floor_elevator2[59]), 
        .out(\eq_47_3/LTV1 [59]) );
  nand2 \eq_47_3/ULTI1_59  ( .a(\eq_47_3/AEQB [59]), .b(\eq_47_3/LTV [59]), 
        .out(\eq_47_3/LTV2 [59]) );
  nand2 \eq_47_3/ULTI2_59  ( .a(\eq_47_3/LTV1 [59]), .b(\eq_47_3/LTV2 [59]), 
        .out(\eq_47_3/LTV [60]) );
  xor2 \eq_47_3/UEQI_60  ( .a(current_floor_output_elevator2[60]), .b(
        destination_floor_elevator2[60]), .out(n2272) );
  nand2 \eq_47_3/UGTI0_60  ( .a(n2271), .b(current_floor_output_elevator2[60]), 
        .out(\eq_47_3/GTV1 [60]) );
  nand2 \eq_47_3/UGTI1_60  ( .a(\eq_47_3/AEQB [60]), .b(\eq_47_3/GTV [60]), 
        .out(\eq_47_3/GTV2 [60]) );
  nand2 \eq_47_3/UGTI2_60  ( .a(\eq_47_3/GTV1 [60]), .b(\eq_47_3/GTV2 [60]), 
        .out(\eq_47_3/GTV [61]) );
  nand2 \eq_47_3/ULTI0_60  ( .a(n2270), .b(destination_floor_elevator2[60]), 
        .out(\eq_47_3/LTV1 [60]) );
  nand2 \eq_47_3/ULTI1_60  ( .a(\eq_47_3/AEQB [60]), .b(\eq_47_3/LTV [60]), 
        .out(\eq_47_3/LTV2 [60]) );
  nand2 \eq_47_3/ULTI2_60  ( .a(\eq_47_3/LTV1 [60]), .b(\eq_47_3/LTV2 [60]), 
        .out(\eq_47_3/LTV [61]) );
  xor2 \eq_47_3/UEQI_61  ( .a(current_floor_output_elevator2[61]), .b(
        destination_floor_elevator2[61]), .out(n2269) );
  nand2 \eq_47_3/UGTI0_61  ( .a(n2268), .b(current_floor_output_elevator2[61]), 
        .out(\eq_47_3/GTV1 [61]) );
  nand2 \eq_47_3/UGTI1_61  ( .a(\eq_47_3/AEQB [61]), .b(\eq_47_3/GTV [61]), 
        .out(\eq_47_3/GTV2 [61]) );
  nand2 \eq_47_3/UGTI2_61  ( .a(\eq_47_3/GTV1 [61]), .b(\eq_47_3/GTV2 [61]), 
        .out(\eq_47_3/GTV [62]) );
  nand2 \eq_47_3/ULTI0_61  ( .a(n2267), .b(destination_floor_elevator2[61]), 
        .out(\eq_47_3/LTV1 [61]) );
  nand2 \eq_47_3/ULTI1_61  ( .a(\eq_47_3/AEQB [61]), .b(\eq_47_3/LTV [61]), 
        .out(\eq_47_3/LTV2 [61]) );
  nand2 \eq_47_3/ULTI2_61  ( .a(\eq_47_3/LTV1 [61]), .b(\eq_47_3/LTV2 [61]), 
        .out(\eq_47_3/LTV [62]) );
  xor2 \eq_47_3/UEQI_62  ( .a(current_floor_output_elevator2[62]), .b(
        destination_floor_elevator2[62]), .out(n2266) );
  nand2 \eq_47_3/UGTI0_62  ( .a(n2265), .b(current_floor_output_elevator2[62]), 
        .out(\eq_47_3/GTV1 [62]) );
  nand2 \eq_47_3/UGTI1_62  ( .a(\eq_47_3/AEQB [62]), .b(\eq_47_3/GTV [62]), 
        .out(\eq_47_3/GTV2 [62]) );
  nand2 \eq_47_3/UGTI2_62  ( .a(\eq_47_3/GTV1 [62]), .b(\eq_47_3/GTV2 [62]), 
        .out(\eq_47_3/GTV [63]) );
  nand2 \eq_47_3/ULTI0_62  ( .a(n2264), .b(destination_floor_elevator2[62]), 
        .out(\eq_47_3/LTV1 [62]) );
  nand2 \eq_47_3/ULTI1_62  ( .a(\eq_47_3/AEQB [62]), .b(\eq_47_3/LTV [62]), 
        .out(\eq_47_3/LTV2 [62]) );
  nand2 \eq_47_3/ULTI2_62  ( .a(\eq_47_3/LTV1 [62]), .b(\eq_47_3/LTV2 [62]), 
        .out(\eq_47_3/LTV [63]) );
  nor2 \ne_47/UEQ  ( .a(\ne_47/GT ), .b(\ne_47/LT ), .out(\ne_47/EQ ) );
  inv \ne_47/UNE  ( .in(\ne_47/EQ ), .out(N15) );
  nand2 \ne_47/UNGT0  ( .a(final_floor_elevator1[0]), .b(n2263), .out(n2262)
         );
  nand2 \ne_47/UNLT0  ( .a(requested_floor[0]), .b(n2261), .out(n2260) );
  xor2 \ne_47/UEQI  ( .a(\ne_47/SA ), .b(\ne_47/SB ), .out(n2259) );
  nand2 \ne_47/UGTI0  ( .a(n2258), .b(\ne_47/SA ), .out(\ne_47/GTV1 [63]) );
  nand2 \ne_47/UGTI1  ( .a(\ne_47/AEQB [63]), .b(\ne_47/GTV [63]), .out(
        \ne_47/GTV2 [63]) );
  nand2 \ne_47/UGTI2  ( .a(\ne_47/GTV1 [63]), .b(\ne_47/GTV2 [63]), .out(
        \ne_47/GT ) );
  nand2 \ne_47/ULTI0  ( .a(n2257), .b(\ne_47/SB ), .out(\ne_47/LTV1 [63]) );
  nand2 \ne_47/ULTI1  ( .a(\ne_47/AEQB [63]), .b(\ne_47/LTV [63]), .out(
        \ne_47/LTV2 [63]) );
  nand2 \ne_47/ULTI2  ( .a(\ne_47/LTV1 [63]), .b(\ne_47/LTV2 [63]), .out(
        \ne_47/LT ) );
  xor2 \ne_47/UEQI_1  ( .a(final_floor_elevator1[1]), .b(requested_floor[1]), 
        .out(n2256) );
  nand2 \ne_47/UGTI0_1  ( .a(n2255), .b(final_floor_elevator1[1]), .out(
        \ne_47/GTV1 [1]) );
  nand2 \ne_47/UGTI1_1  ( .a(\ne_47/AEQB [1]), .b(\ne_47/GTV [1]), .out(
        \ne_47/GTV2 [1]) );
  nand2 \ne_47/UGTI2_1  ( .a(\ne_47/GTV1 [1]), .b(\ne_47/GTV2 [1]), .out(
        \ne_47/GTV [2]) );
  nand2 \ne_47/ULTI0_1  ( .a(n2254), .b(requested_floor[1]), .out(
        \ne_47/LTV1 [1]) );
  nand2 \ne_47/ULTI1_1  ( .a(\ne_47/AEQB [1]), .b(\ne_47/LTV [1]), .out(
        \ne_47/LTV2 [1]) );
  nand2 \ne_47/ULTI2_1  ( .a(\ne_47/LTV1 [1]), .b(\ne_47/LTV2 [1]), .out(
        \ne_47/LTV [2]) );
  xor2 \ne_47/UEQI_2  ( .a(final_floor_elevator1[2]), .b(requested_floor[2]), 
        .out(n2253) );
  nand2 \ne_47/UGTI0_2  ( .a(n2252), .b(final_floor_elevator1[2]), .out(
        \ne_47/GTV1 [2]) );
  nand2 \ne_47/UGTI1_2  ( .a(\ne_47/AEQB [2]), .b(\ne_47/GTV [2]), .out(
        \ne_47/GTV2 [2]) );
  nand2 \ne_47/UGTI2_2  ( .a(\ne_47/GTV1 [2]), .b(\ne_47/GTV2 [2]), .out(
        \ne_47/GTV [3]) );
  nand2 \ne_47/ULTI0_2  ( .a(n2251), .b(requested_floor[2]), .out(
        \ne_47/LTV1 [2]) );
  nand2 \ne_47/ULTI1_2  ( .a(\ne_47/AEQB [2]), .b(\ne_47/LTV [2]), .out(
        \ne_47/LTV2 [2]) );
  nand2 \ne_47/ULTI2_2  ( .a(\ne_47/LTV1 [2]), .b(\ne_47/LTV2 [2]), .out(
        \ne_47/LTV [3]) );
  xor2 \ne_47/UEQI_3  ( .a(final_floor_elevator1[3]), .b(requested_floor[3]), 
        .out(n2250) );
  nand2 \ne_47/UGTI0_3  ( .a(n2249), .b(final_floor_elevator1[3]), .out(
        \ne_47/GTV1 [3]) );
  nand2 \ne_47/UGTI1_3  ( .a(\ne_47/AEQB [3]), .b(\ne_47/GTV [3]), .out(
        \ne_47/GTV2 [3]) );
  nand2 \ne_47/UGTI2_3  ( .a(\ne_47/GTV1 [3]), .b(\ne_47/GTV2 [3]), .out(
        \ne_47/GTV [4]) );
  nand2 \ne_47/ULTI0_3  ( .a(n2248), .b(requested_floor[3]), .out(
        \ne_47/LTV1 [3]) );
  nand2 \ne_47/ULTI1_3  ( .a(\ne_47/AEQB [3]), .b(\ne_47/LTV [3]), .out(
        \ne_47/LTV2 [3]) );
  nand2 \ne_47/ULTI2_3  ( .a(\ne_47/LTV1 [3]), .b(\ne_47/LTV2 [3]), .out(
        \ne_47/LTV [4]) );
  xor2 \ne_47/UEQI_4  ( .a(final_floor_elevator1[4]), .b(requested_floor[4]), 
        .out(n2247) );
  nand2 \ne_47/UGTI0_4  ( .a(n2246), .b(final_floor_elevator1[4]), .out(
        \ne_47/GTV1 [4]) );
  nand2 \ne_47/UGTI1_4  ( .a(\ne_47/AEQB [4]), .b(\ne_47/GTV [4]), .out(
        \ne_47/GTV2 [4]) );
  nand2 \ne_47/UGTI2_4  ( .a(\ne_47/GTV1 [4]), .b(\ne_47/GTV2 [4]), .out(
        \ne_47/GTV [5]) );
  nand2 \ne_47/ULTI0_4  ( .a(n2245), .b(requested_floor[4]), .out(
        \ne_47/LTV1 [4]) );
  nand2 \ne_47/ULTI1_4  ( .a(\ne_47/AEQB [4]), .b(\ne_47/LTV [4]), .out(
        \ne_47/LTV2 [4]) );
  nand2 \ne_47/ULTI2_4  ( .a(\ne_47/LTV1 [4]), .b(\ne_47/LTV2 [4]), .out(
        \ne_47/LTV [5]) );
  xor2 \ne_47/UEQI_5  ( .a(final_floor_elevator1[5]), .b(requested_floor[5]), 
        .out(n2244) );
  nand2 \ne_47/UGTI0_5  ( .a(n2243), .b(final_floor_elevator1[5]), .out(
        \ne_47/GTV1 [5]) );
  nand2 \ne_47/UGTI1_5  ( .a(\ne_47/AEQB [5]), .b(\ne_47/GTV [5]), .out(
        \ne_47/GTV2 [5]) );
  nand2 \ne_47/UGTI2_5  ( .a(\ne_47/GTV1 [5]), .b(\ne_47/GTV2 [5]), .out(
        \ne_47/GTV [6]) );
  nand2 \ne_47/ULTI0_5  ( .a(n2242), .b(requested_floor[5]), .out(
        \ne_47/LTV1 [5]) );
  nand2 \ne_47/ULTI1_5  ( .a(\ne_47/AEQB [5]), .b(\ne_47/LTV [5]), .out(
        \ne_47/LTV2 [5]) );
  nand2 \ne_47/ULTI2_5  ( .a(\ne_47/LTV1 [5]), .b(\ne_47/LTV2 [5]), .out(
        \ne_47/LTV [6]) );
  xor2 \ne_47/UEQI_6  ( .a(final_floor_elevator1[6]), .b(requested_floor[6]), 
        .out(n2241) );
  nand2 \ne_47/UGTI0_6  ( .a(n2240), .b(final_floor_elevator1[6]), .out(
        \ne_47/GTV1 [6]) );
  nand2 \ne_47/UGTI1_6  ( .a(\ne_47/AEQB [6]), .b(\ne_47/GTV [6]), .out(
        \ne_47/GTV2 [6]) );
  nand2 \ne_47/UGTI2_6  ( .a(\ne_47/GTV1 [6]), .b(\ne_47/GTV2 [6]), .out(
        \ne_47/GTV [7]) );
  nand2 \ne_47/ULTI0_6  ( .a(n2239), .b(requested_floor[6]), .out(
        \ne_47/LTV1 [6]) );
  nand2 \ne_47/ULTI1_6  ( .a(\ne_47/AEQB [6]), .b(\ne_47/LTV [6]), .out(
        \ne_47/LTV2 [6]) );
  nand2 \ne_47/ULTI2_6  ( .a(\ne_47/LTV1 [6]), .b(\ne_47/LTV2 [6]), .out(
        \ne_47/LTV [7]) );
  xor2 \ne_47/UEQI_7  ( .a(final_floor_elevator1[7]), .b(requested_floor[7]), 
        .out(n2238) );
  nand2 \ne_47/UGTI0_7  ( .a(n2237), .b(final_floor_elevator1[7]), .out(
        \ne_47/GTV1 [7]) );
  nand2 \ne_47/UGTI1_7  ( .a(\ne_47/AEQB [7]), .b(\ne_47/GTV [7]), .out(
        \ne_47/GTV2 [7]) );
  nand2 \ne_47/UGTI2_7  ( .a(\ne_47/GTV1 [7]), .b(\ne_47/GTV2 [7]), .out(
        \ne_47/GTV [8]) );
  nand2 \ne_47/ULTI0_7  ( .a(n2236), .b(requested_floor[7]), .out(
        \ne_47/LTV1 [7]) );
  nand2 \ne_47/ULTI1_7  ( .a(\ne_47/AEQB [7]), .b(\ne_47/LTV [7]), .out(
        \ne_47/LTV2 [7]) );
  nand2 \ne_47/ULTI2_7  ( .a(\ne_47/LTV1 [7]), .b(\ne_47/LTV2 [7]), .out(
        \ne_47/LTV [8]) );
  xor2 \ne_47/UEQI_8  ( .a(final_floor_elevator1[8]), .b(requested_floor[8]), 
        .out(n2235) );
  nand2 \ne_47/UGTI0_8  ( .a(n2234), .b(final_floor_elevator1[8]), .out(
        \ne_47/GTV1 [8]) );
  nand2 \ne_47/UGTI1_8  ( .a(\ne_47/AEQB [8]), .b(\ne_47/GTV [8]), .out(
        \ne_47/GTV2 [8]) );
  nand2 \ne_47/UGTI2_8  ( .a(\ne_47/GTV1 [8]), .b(\ne_47/GTV2 [8]), .out(
        \ne_47/GTV [9]) );
  nand2 \ne_47/ULTI0_8  ( .a(n2233), .b(requested_floor[8]), .out(
        \ne_47/LTV1 [8]) );
  nand2 \ne_47/ULTI1_8  ( .a(\ne_47/AEQB [8]), .b(\ne_47/LTV [8]), .out(
        \ne_47/LTV2 [8]) );
  nand2 \ne_47/ULTI2_8  ( .a(\ne_47/LTV1 [8]), .b(\ne_47/LTV2 [8]), .out(
        \ne_47/LTV [9]) );
  xor2 \ne_47/UEQI_9  ( .a(final_floor_elevator1[9]), .b(requested_floor[9]), 
        .out(n2232) );
  nand2 \ne_47/UGTI0_9  ( .a(n2231), .b(final_floor_elevator1[9]), .out(
        \ne_47/GTV1 [9]) );
  nand2 \ne_47/UGTI1_9  ( .a(\ne_47/AEQB [9]), .b(\ne_47/GTV [9]), .out(
        \ne_47/GTV2 [9]) );
  nand2 \ne_47/UGTI2_9  ( .a(\ne_47/GTV1 [9]), .b(\ne_47/GTV2 [9]), .out(
        \ne_47/GTV [10]) );
  nand2 \ne_47/ULTI0_9  ( .a(n2230), .b(requested_floor[9]), .out(
        \ne_47/LTV1 [9]) );
  nand2 \ne_47/ULTI1_9  ( .a(\ne_47/AEQB [9]), .b(\ne_47/LTV [9]), .out(
        \ne_47/LTV2 [9]) );
  nand2 \ne_47/ULTI2_9  ( .a(\ne_47/LTV1 [9]), .b(\ne_47/LTV2 [9]), .out(
        \ne_47/LTV [10]) );
  xor2 \ne_47/UEQI_10  ( .a(final_floor_elevator1[10]), .b(requested_floor[10]), .out(n2229) );
  nand2 \ne_47/UGTI0_10  ( .a(n2228), .b(final_floor_elevator1[10]), .out(
        \ne_47/GTV1 [10]) );
  nand2 \ne_47/UGTI1_10  ( .a(\ne_47/AEQB [10]), .b(\ne_47/GTV [10]), .out(
        \ne_47/GTV2 [10]) );
  nand2 \ne_47/UGTI2_10  ( .a(\ne_47/GTV1 [10]), .b(\ne_47/GTV2 [10]), .out(
        \ne_47/GTV [11]) );
  nand2 \ne_47/ULTI0_10  ( .a(n2227), .b(requested_floor[10]), .out(
        \ne_47/LTV1 [10]) );
  nand2 \ne_47/ULTI1_10  ( .a(\ne_47/AEQB [10]), .b(\ne_47/LTV [10]), .out(
        \ne_47/LTV2 [10]) );
  nand2 \ne_47/ULTI2_10  ( .a(\ne_47/LTV1 [10]), .b(\ne_47/LTV2 [10]), .out(
        \ne_47/LTV [11]) );
  xor2 \ne_47/UEQI_11  ( .a(final_floor_elevator1[11]), .b(requested_floor[11]), .out(n2226) );
  nand2 \ne_47/UGTI0_11  ( .a(n2225), .b(final_floor_elevator1[11]), .out(
        \ne_47/GTV1 [11]) );
  nand2 \ne_47/UGTI1_11  ( .a(\ne_47/AEQB [11]), .b(\ne_47/GTV [11]), .out(
        \ne_47/GTV2 [11]) );
  nand2 \ne_47/UGTI2_11  ( .a(\ne_47/GTV1 [11]), .b(\ne_47/GTV2 [11]), .out(
        \ne_47/GTV [12]) );
  nand2 \ne_47/ULTI0_11  ( .a(n2224), .b(requested_floor[11]), .out(
        \ne_47/LTV1 [11]) );
  nand2 \ne_47/ULTI1_11  ( .a(\ne_47/AEQB [11]), .b(\ne_47/LTV [11]), .out(
        \ne_47/LTV2 [11]) );
  nand2 \ne_47/ULTI2_11  ( .a(\ne_47/LTV1 [11]), .b(\ne_47/LTV2 [11]), .out(
        \ne_47/LTV [12]) );
  xor2 \ne_47/UEQI_12  ( .a(final_floor_elevator1[12]), .b(requested_floor[12]), .out(n2223) );
  nand2 \ne_47/UGTI0_12  ( .a(n2222), .b(final_floor_elevator1[12]), .out(
        \ne_47/GTV1 [12]) );
  nand2 \ne_47/UGTI1_12  ( .a(\ne_47/AEQB [12]), .b(\ne_47/GTV [12]), .out(
        \ne_47/GTV2 [12]) );
  nand2 \ne_47/UGTI2_12  ( .a(\ne_47/GTV1 [12]), .b(\ne_47/GTV2 [12]), .out(
        \ne_47/GTV [13]) );
  nand2 \ne_47/ULTI0_12  ( .a(n2221), .b(requested_floor[12]), .out(
        \ne_47/LTV1 [12]) );
  nand2 \ne_47/ULTI1_12  ( .a(\ne_47/AEQB [12]), .b(\ne_47/LTV [12]), .out(
        \ne_47/LTV2 [12]) );
  nand2 \ne_47/ULTI2_12  ( .a(\ne_47/LTV1 [12]), .b(\ne_47/LTV2 [12]), .out(
        \ne_47/LTV [13]) );
  xor2 \ne_47/UEQI_13  ( .a(final_floor_elevator1[13]), .b(requested_floor[13]), .out(n2220) );
  nand2 \ne_47/UGTI0_13  ( .a(n2219), .b(final_floor_elevator1[13]), .out(
        \ne_47/GTV1 [13]) );
  nand2 \ne_47/UGTI1_13  ( .a(\ne_47/AEQB [13]), .b(\ne_47/GTV [13]), .out(
        \ne_47/GTV2 [13]) );
  nand2 \ne_47/UGTI2_13  ( .a(\ne_47/GTV1 [13]), .b(\ne_47/GTV2 [13]), .out(
        \ne_47/GTV [14]) );
  nand2 \ne_47/ULTI0_13  ( .a(n2218), .b(requested_floor[13]), .out(
        \ne_47/LTV1 [13]) );
  nand2 \ne_47/ULTI1_13  ( .a(\ne_47/AEQB [13]), .b(\ne_47/LTV [13]), .out(
        \ne_47/LTV2 [13]) );
  nand2 \ne_47/ULTI2_13  ( .a(\ne_47/LTV1 [13]), .b(\ne_47/LTV2 [13]), .out(
        \ne_47/LTV [14]) );
  xor2 \ne_47/UEQI_14  ( .a(final_floor_elevator1[14]), .b(requested_floor[14]), .out(n2217) );
  nand2 \ne_47/UGTI0_14  ( .a(n2216), .b(final_floor_elevator1[14]), .out(
        \ne_47/GTV1 [14]) );
  nand2 \ne_47/UGTI1_14  ( .a(\ne_47/AEQB [14]), .b(\ne_47/GTV [14]), .out(
        \ne_47/GTV2 [14]) );
  nand2 \ne_47/UGTI2_14  ( .a(\ne_47/GTV1 [14]), .b(\ne_47/GTV2 [14]), .out(
        \ne_47/GTV [15]) );
  nand2 \ne_47/ULTI0_14  ( .a(n2215), .b(requested_floor[14]), .out(
        \ne_47/LTV1 [14]) );
  nand2 \ne_47/ULTI1_14  ( .a(\ne_47/AEQB [14]), .b(\ne_47/LTV [14]), .out(
        \ne_47/LTV2 [14]) );
  nand2 \ne_47/ULTI2_14  ( .a(\ne_47/LTV1 [14]), .b(\ne_47/LTV2 [14]), .out(
        \ne_47/LTV [15]) );
  xor2 \ne_47/UEQI_15  ( .a(final_floor_elevator1[15]), .b(requested_floor[15]), .out(n2214) );
  nand2 \ne_47/UGTI0_15  ( .a(n2213), .b(final_floor_elevator1[15]), .out(
        \ne_47/GTV1 [15]) );
  nand2 \ne_47/UGTI1_15  ( .a(\ne_47/AEQB [15]), .b(\ne_47/GTV [15]), .out(
        \ne_47/GTV2 [15]) );
  nand2 \ne_47/UGTI2_15  ( .a(\ne_47/GTV1 [15]), .b(\ne_47/GTV2 [15]), .out(
        \ne_47/GTV [16]) );
  nand2 \ne_47/ULTI0_15  ( .a(n2212), .b(requested_floor[15]), .out(
        \ne_47/LTV1 [15]) );
  nand2 \ne_47/ULTI1_15  ( .a(\ne_47/AEQB [15]), .b(\ne_47/LTV [15]), .out(
        \ne_47/LTV2 [15]) );
  nand2 \ne_47/ULTI2_15  ( .a(\ne_47/LTV1 [15]), .b(\ne_47/LTV2 [15]), .out(
        \ne_47/LTV [16]) );
  xor2 \ne_47/UEQI_16  ( .a(final_floor_elevator1[16]), .b(requested_floor[16]), .out(n2211) );
  nand2 \ne_47/UGTI0_16  ( .a(n2210), .b(final_floor_elevator1[16]), .out(
        \ne_47/GTV1 [16]) );
  nand2 \ne_47/UGTI1_16  ( .a(\ne_47/AEQB [16]), .b(\ne_47/GTV [16]), .out(
        \ne_47/GTV2 [16]) );
  nand2 \ne_47/UGTI2_16  ( .a(\ne_47/GTV1 [16]), .b(\ne_47/GTV2 [16]), .out(
        \ne_47/GTV [17]) );
  nand2 \ne_47/ULTI0_16  ( .a(n2209), .b(requested_floor[16]), .out(
        \ne_47/LTV1 [16]) );
  nand2 \ne_47/ULTI1_16  ( .a(\ne_47/AEQB [16]), .b(\ne_47/LTV [16]), .out(
        \ne_47/LTV2 [16]) );
  nand2 \ne_47/ULTI2_16  ( .a(\ne_47/LTV1 [16]), .b(\ne_47/LTV2 [16]), .out(
        \ne_47/LTV [17]) );
  xor2 \ne_47/UEQI_17  ( .a(final_floor_elevator1[17]), .b(requested_floor[17]), .out(n2208) );
  nand2 \ne_47/UGTI0_17  ( .a(n2207), .b(final_floor_elevator1[17]), .out(
        \ne_47/GTV1 [17]) );
  nand2 \ne_47/UGTI1_17  ( .a(\ne_47/AEQB [17]), .b(\ne_47/GTV [17]), .out(
        \ne_47/GTV2 [17]) );
  nand2 \ne_47/UGTI2_17  ( .a(\ne_47/GTV1 [17]), .b(\ne_47/GTV2 [17]), .out(
        \ne_47/GTV [18]) );
  nand2 \ne_47/ULTI0_17  ( .a(n2206), .b(requested_floor[17]), .out(
        \ne_47/LTV1 [17]) );
  nand2 \ne_47/ULTI1_17  ( .a(\ne_47/AEQB [17]), .b(\ne_47/LTV [17]), .out(
        \ne_47/LTV2 [17]) );
  nand2 \ne_47/ULTI2_17  ( .a(\ne_47/LTV1 [17]), .b(\ne_47/LTV2 [17]), .out(
        \ne_47/LTV [18]) );
  xor2 \ne_47/UEQI_18  ( .a(final_floor_elevator1[18]), .b(requested_floor[18]), .out(n2205) );
  nand2 \ne_47/UGTI0_18  ( .a(n2204), .b(final_floor_elevator1[18]), .out(
        \ne_47/GTV1 [18]) );
  nand2 \ne_47/UGTI1_18  ( .a(\ne_47/AEQB [18]), .b(\ne_47/GTV [18]), .out(
        \ne_47/GTV2 [18]) );
  nand2 \ne_47/UGTI2_18  ( .a(\ne_47/GTV1 [18]), .b(\ne_47/GTV2 [18]), .out(
        \ne_47/GTV [19]) );
  nand2 \ne_47/ULTI0_18  ( .a(n2203), .b(requested_floor[18]), .out(
        \ne_47/LTV1 [18]) );
  nand2 \ne_47/ULTI1_18  ( .a(\ne_47/AEQB [18]), .b(\ne_47/LTV [18]), .out(
        \ne_47/LTV2 [18]) );
  nand2 \ne_47/ULTI2_18  ( .a(\ne_47/LTV1 [18]), .b(\ne_47/LTV2 [18]), .out(
        \ne_47/LTV [19]) );
  xor2 \ne_47/UEQI_19  ( .a(final_floor_elevator1[19]), .b(requested_floor[19]), .out(n2202) );
  nand2 \ne_47/UGTI0_19  ( .a(n2201), .b(final_floor_elevator1[19]), .out(
        \ne_47/GTV1 [19]) );
  nand2 \ne_47/UGTI1_19  ( .a(\ne_47/AEQB [19]), .b(\ne_47/GTV [19]), .out(
        \ne_47/GTV2 [19]) );
  nand2 \ne_47/UGTI2_19  ( .a(\ne_47/GTV1 [19]), .b(\ne_47/GTV2 [19]), .out(
        \ne_47/GTV [20]) );
  nand2 \ne_47/ULTI0_19  ( .a(n2200), .b(requested_floor[19]), .out(
        \ne_47/LTV1 [19]) );
  nand2 \ne_47/ULTI1_19  ( .a(\ne_47/AEQB [19]), .b(\ne_47/LTV [19]), .out(
        \ne_47/LTV2 [19]) );
  nand2 \ne_47/ULTI2_19  ( .a(\ne_47/LTV1 [19]), .b(\ne_47/LTV2 [19]), .out(
        \ne_47/LTV [20]) );
  xor2 \ne_47/UEQI_20  ( .a(final_floor_elevator1[20]), .b(requested_floor[20]), .out(n2199) );
  nand2 \ne_47/UGTI0_20  ( .a(n2198), .b(final_floor_elevator1[20]), .out(
        \ne_47/GTV1 [20]) );
  nand2 \ne_47/UGTI1_20  ( .a(\ne_47/AEQB [20]), .b(\ne_47/GTV [20]), .out(
        \ne_47/GTV2 [20]) );
  nand2 \ne_47/UGTI2_20  ( .a(\ne_47/GTV1 [20]), .b(\ne_47/GTV2 [20]), .out(
        \ne_47/GTV [21]) );
  nand2 \ne_47/ULTI0_20  ( .a(n2197), .b(requested_floor[20]), .out(
        \ne_47/LTV1 [20]) );
  nand2 \ne_47/ULTI1_20  ( .a(\ne_47/AEQB [20]), .b(\ne_47/LTV [20]), .out(
        \ne_47/LTV2 [20]) );
  nand2 \ne_47/ULTI2_20  ( .a(\ne_47/LTV1 [20]), .b(\ne_47/LTV2 [20]), .out(
        \ne_47/LTV [21]) );
  xor2 \ne_47/UEQI_21  ( .a(final_floor_elevator1[21]), .b(requested_floor[21]), .out(n2196) );
  nand2 \ne_47/UGTI0_21  ( .a(n2195), .b(final_floor_elevator1[21]), .out(
        \ne_47/GTV1 [21]) );
  nand2 \ne_47/UGTI1_21  ( .a(\ne_47/AEQB [21]), .b(\ne_47/GTV [21]), .out(
        \ne_47/GTV2 [21]) );
  nand2 \ne_47/UGTI2_21  ( .a(\ne_47/GTV1 [21]), .b(\ne_47/GTV2 [21]), .out(
        \ne_47/GTV [22]) );
  nand2 \ne_47/ULTI0_21  ( .a(n2194), .b(requested_floor[21]), .out(
        \ne_47/LTV1 [21]) );
  nand2 \ne_47/ULTI1_21  ( .a(\ne_47/AEQB [21]), .b(\ne_47/LTV [21]), .out(
        \ne_47/LTV2 [21]) );
  nand2 \ne_47/ULTI2_21  ( .a(\ne_47/LTV1 [21]), .b(\ne_47/LTV2 [21]), .out(
        \ne_47/LTV [22]) );
  xor2 \ne_47/UEQI_22  ( .a(final_floor_elevator1[22]), .b(requested_floor[22]), .out(n2193) );
  nand2 \ne_47/UGTI0_22  ( .a(n2192), .b(final_floor_elevator1[22]), .out(
        \ne_47/GTV1 [22]) );
  nand2 \ne_47/UGTI1_22  ( .a(\ne_47/AEQB [22]), .b(\ne_47/GTV [22]), .out(
        \ne_47/GTV2 [22]) );
  nand2 \ne_47/UGTI2_22  ( .a(\ne_47/GTV1 [22]), .b(\ne_47/GTV2 [22]), .out(
        \ne_47/GTV [23]) );
  nand2 \ne_47/ULTI0_22  ( .a(n2191), .b(requested_floor[22]), .out(
        \ne_47/LTV1 [22]) );
  nand2 \ne_47/ULTI1_22  ( .a(\ne_47/AEQB [22]), .b(\ne_47/LTV [22]), .out(
        \ne_47/LTV2 [22]) );
  nand2 \ne_47/ULTI2_22  ( .a(\ne_47/LTV1 [22]), .b(\ne_47/LTV2 [22]), .out(
        \ne_47/LTV [23]) );
  xor2 \ne_47/UEQI_23  ( .a(final_floor_elevator1[23]), .b(requested_floor[23]), .out(n2190) );
  nand2 \ne_47/UGTI0_23  ( .a(n2189), .b(final_floor_elevator1[23]), .out(
        \ne_47/GTV1 [23]) );
  nand2 \ne_47/UGTI1_23  ( .a(\ne_47/AEQB [23]), .b(\ne_47/GTV [23]), .out(
        \ne_47/GTV2 [23]) );
  nand2 \ne_47/UGTI2_23  ( .a(\ne_47/GTV1 [23]), .b(\ne_47/GTV2 [23]), .out(
        \ne_47/GTV [24]) );
  nand2 \ne_47/ULTI0_23  ( .a(n2188), .b(requested_floor[23]), .out(
        \ne_47/LTV1 [23]) );
  nand2 \ne_47/ULTI1_23  ( .a(\ne_47/AEQB [23]), .b(\ne_47/LTV [23]), .out(
        \ne_47/LTV2 [23]) );
  nand2 \ne_47/ULTI2_23  ( .a(\ne_47/LTV1 [23]), .b(\ne_47/LTV2 [23]), .out(
        \ne_47/LTV [24]) );
  xor2 \ne_47/UEQI_24  ( .a(final_floor_elevator1[24]), .b(requested_floor[24]), .out(n2187) );
  nand2 \ne_47/UGTI0_24  ( .a(n2186), .b(final_floor_elevator1[24]), .out(
        \ne_47/GTV1 [24]) );
  nand2 \ne_47/UGTI1_24  ( .a(\ne_47/AEQB [24]), .b(\ne_47/GTV [24]), .out(
        \ne_47/GTV2 [24]) );
  nand2 \ne_47/UGTI2_24  ( .a(\ne_47/GTV1 [24]), .b(\ne_47/GTV2 [24]), .out(
        \ne_47/GTV [25]) );
  nand2 \ne_47/ULTI0_24  ( .a(n2185), .b(requested_floor[24]), .out(
        \ne_47/LTV1 [24]) );
  nand2 \ne_47/ULTI1_24  ( .a(\ne_47/AEQB [24]), .b(\ne_47/LTV [24]), .out(
        \ne_47/LTV2 [24]) );
  nand2 \ne_47/ULTI2_24  ( .a(\ne_47/LTV1 [24]), .b(\ne_47/LTV2 [24]), .out(
        \ne_47/LTV [25]) );
  xor2 \ne_47/UEQI_25  ( .a(final_floor_elevator1[25]), .b(requested_floor[25]), .out(n2184) );
  nand2 \ne_47/UGTI0_25  ( .a(n2183), .b(final_floor_elevator1[25]), .out(
        \ne_47/GTV1 [25]) );
  nand2 \ne_47/UGTI1_25  ( .a(\ne_47/AEQB [25]), .b(\ne_47/GTV [25]), .out(
        \ne_47/GTV2 [25]) );
  nand2 \ne_47/UGTI2_25  ( .a(\ne_47/GTV1 [25]), .b(\ne_47/GTV2 [25]), .out(
        \ne_47/GTV [26]) );
  nand2 \ne_47/ULTI0_25  ( .a(n2182), .b(requested_floor[25]), .out(
        \ne_47/LTV1 [25]) );
  nand2 \ne_47/ULTI1_25  ( .a(\ne_47/AEQB [25]), .b(\ne_47/LTV [25]), .out(
        \ne_47/LTV2 [25]) );
  nand2 \ne_47/ULTI2_25  ( .a(\ne_47/LTV1 [25]), .b(\ne_47/LTV2 [25]), .out(
        \ne_47/LTV [26]) );
  xor2 \ne_47/UEQI_26  ( .a(final_floor_elevator1[26]), .b(requested_floor[26]), .out(n2181) );
  nand2 \ne_47/UGTI0_26  ( .a(n2180), .b(final_floor_elevator1[26]), .out(
        \ne_47/GTV1 [26]) );
  nand2 \ne_47/UGTI1_26  ( .a(\ne_47/AEQB [26]), .b(\ne_47/GTV [26]), .out(
        \ne_47/GTV2 [26]) );
  nand2 \ne_47/UGTI2_26  ( .a(\ne_47/GTV1 [26]), .b(\ne_47/GTV2 [26]), .out(
        \ne_47/GTV [27]) );
  nand2 \ne_47/ULTI0_26  ( .a(n2179), .b(requested_floor[26]), .out(
        \ne_47/LTV1 [26]) );
  nand2 \ne_47/ULTI1_26  ( .a(\ne_47/AEQB [26]), .b(\ne_47/LTV [26]), .out(
        \ne_47/LTV2 [26]) );
  nand2 \ne_47/ULTI2_26  ( .a(\ne_47/LTV1 [26]), .b(\ne_47/LTV2 [26]), .out(
        \ne_47/LTV [27]) );
  xor2 \ne_47/UEQI_27  ( .a(final_floor_elevator1[27]), .b(requested_floor[27]), .out(n2178) );
  nand2 \ne_47/UGTI0_27  ( .a(n2177), .b(final_floor_elevator1[27]), .out(
        \ne_47/GTV1 [27]) );
  nand2 \ne_47/UGTI1_27  ( .a(\ne_47/AEQB [27]), .b(\ne_47/GTV [27]), .out(
        \ne_47/GTV2 [27]) );
  nand2 \ne_47/UGTI2_27  ( .a(\ne_47/GTV1 [27]), .b(\ne_47/GTV2 [27]), .out(
        \ne_47/GTV [28]) );
  nand2 \ne_47/ULTI0_27  ( .a(n2176), .b(requested_floor[27]), .out(
        \ne_47/LTV1 [27]) );
  nand2 \ne_47/ULTI1_27  ( .a(\ne_47/AEQB [27]), .b(\ne_47/LTV [27]), .out(
        \ne_47/LTV2 [27]) );
  nand2 \ne_47/ULTI2_27  ( .a(\ne_47/LTV1 [27]), .b(\ne_47/LTV2 [27]), .out(
        \ne_47/LTV [28]) );
  xor2 \ne_47/UEQI_28  ( .a(final_floor_elevator1[28]), .b(requested_floor[28]), .out(n2175) );
  nand2 \ne_47/UGTI0_28  ( .a(n2174), .b(final_floor_elevator1[28]), .out(
        \ne_47/GTV1 [28]) );
  nand2 \ne_47/UGTI1_28  ( .a(\ne_47/AEQB [28]), .b(\ne_47/GTV [28]), .out(
        \ne_47/GTV2 [28]) );
  nand2 \ne_47/UGTI2_28  ( .a(\ne_47/GTV1 [28]), .b(\ne_47/GTV2 [28]), .out(
        \ne_47/GTV [29]) );
  nand2 \ne_47/ULTI0_28  ( .a(n2173), .b(requested_floor[28]), .out(
        \ne_47/LTV1 [28]) );
  nand2 \ne_47/ULTI1_28  ( .a(\ne_47/AEQB [28]), .b(\ne_47/LTV [28]), .out(
        \ne_47/LTV2 [28]) );
  nand2 \ne_47/ULTI2_28  ( .a(\ne_47/LTV1 [28]), .b(\ne_47/LTV2 [28]), .out(
        \ne_47/LTV [29]) );
  xor2 \ne_47/UEQI_29  ( .a(final_floor_elevator1[29]), .b(requested_floor[29]), .out(n2172) );
  nand2 \ne_47/UGTI0_29  ( .a(n2171), .b(final_floor_elevator1[29]), .out(
        \ne_47/GTV1 [29]) );
  nand2 \ne_47/UGTI1_29  ( .a(\ne_47/AEQB [29]), .b(\ne_47/GTV [29]), .out(
        \ne_47/GTV2 [29]) );
  nand2 \ne_47/UGTI2_29  ( .a(\ne_47/GTV1 [29]), .b(\ne_47/GTV2 [29]), .out(
        \ne_47/GTV [30]) );
  nand2 \ne_47/ULTI0_29  ( .a(n2170), .b(requested_floor[29]), .out(
        \ne_47/LTV1 [29]) );
  nand2 \ne_47/ULTI1_29  ( .a(\ne_47/AEQB [29]), .b(\ne_47/LTV [29]), .out(
        \ne_47/LTV2 [29]) );
  nand2 \ne_47/ULTI2_29  ( .a(\ne_47/LTV1 [29]), .b(\ne_47/LTV2 [29]), .out(
        \ne_47/LTV [30]) );
  xor2 \ne_47/UEQI_30  ( .a(final_floor_elevator1[30]), .b(requested_floor[30]), .out(n2169) );
  nand2 \ne_47/UGTI0_30  ( .a(n2168), .b(final_floor_elevator1[30]), .out(
        \ne_47/GTV1 [30]) );
  nand2 \ne_47/UGTI1_30  ( .a(\ne_47/AEQB [30]), .b(\ne_47/GTV [30]), .out(
        \ne_47/GTV2 [30]) );
  nand2 \ne_47/UGTI2_30  ( .a(\ne_47/GTV1 [30]), .b(\ne_47/GTV2 [30]), .out(
        \ne_47/GTV [31]) );
  nand2 \ne_47/ULTI0_30  ( .a(n2167), .b(requested_floor[30]), .out(
        \ne_47/LTV1 [30]) );
  nand2 \ne_47/ULTI1_30  ( .a(\ne_47/AEQB [30]), .b(\ne_47/LTV [30]), .out(
        \ne_47/LTV2 [30]) );
  nand2 \ne_47/ULTI2_30  ( .a(\ne_47/LTV1 [30]), .b(\ne_47/LTV2 [30]), .out(
        \ne_47/LTV [31]) );
  xor2 \ne_47/UEQI_31  ( .a(final_floor_elevator1[31]), .b(requested_floor[31]), .out(n2166) );
  nand2 \ne_47/UGTI0_31  ( .a(n2165), .b(final_floor_elevator1[31]), .out(
        \ne_47/GTV1 [31]) );
  nand2 \ne_47/UGTI1_31  ( .a(\ne_47/AEQB [31]), .b(\ne_47/GTV [31]), .out(
        \ne_47/GTV2 [31]) );
  nand2 \ne_47/UGTI2_31  ( .a(\ne_47/GTV1 [31]), .b(\ne_47/GTV2 [31]), .out(
        \ne_47/GTV [32]) );
  nand2 \ne_47/ULTI0_31  ( .a(n2164), .b(requested_floor[31]), .out(
        \ne_47/LTV1 [31]) );
  nand2 \ne_47/ULTI1_31  ( .a(\ne_47/AEQB [31]), .b(\ne_47/LTV [31]), .out(
        \ne_47/LTV2 [31]) );
  nand2 \ne_47/ULTI2_31  ( .a(\ne_47/LTV1 [31]), .b(\ne_47/LTV2 [31]), .out(
        \ne_47/LTV [32]) );
  xor2 \ne_47/UEQI_32  ( .a(final_floor_elevator1[32]), .b(requested_floor[32]), .out(n2163) );
  nand2 \ne_47/UGTI0_32  ( .a(n2162), .b(final_floor_elevator1[32]), .out(
        \ne_47/GTV1 [32]) );
  nand2 \ne_47/UGTI1_32  ( .a(\ne_47/AEQB [32]), .b(\ne_47/GTV [32]), .out(
        \ne_47/GTV2 [32]) );
  nand2 \ne_47/UGTI2_32  ( .a(\ne_47/GTV1 [32]), .b(\ne_47/GTV2 [32]), .out(
        \ne_47/GTV [33]) );
  nand2 \ne_47/ULTI0_32  ( .a(n2161), .b(requested_floor[32]), .out(
        \ne_47/LTV1 [32]) );
  nand2 \ne_47/ULTI1_32  ( .a(\ne_47/AEQB [32]), .b(\ne_47/LTV [32]), .out(
        \ne_47/LTV2 [32]) );
  nand2 \ne_47/ULTI2_32  ( .a(\ne_47/LTV1 [32]), .b(\ne_47/LTV2 [32]), .out(
        \ne_47/LTV [33]) );
  xor2 \ne_47/UEQI_33  ( .a(final_floor_elevator1[33]), .b(requested_floor[33]), .out(n2160) );
  nand2 \ne_47/UGTI0_33  ( .a(n2159), .b(final_floor_elevator1[33]), .out(
        \ne_47/GTV1 [33]) );
  nand2 \ne_47/UGTI1_33  ( .a(\ne_47/AEQB [33]), .b(\ne_47/GTV [33]), .out(
        \ne_47/GTV2 [33]) );
  nand2 \ne_47/UGTI2_33  ( .a(\ne_47/GTV1 [33]), .b(\ne_47/GTV2 [33]), .out(
        \ne_47/GTV [34]) );
  nand2 \ne_47/ULTI0_33  ( .a(n2158), .b(requested_floor[33]), .out(
        \ne_47/LTV1 [33]) );
  nand2 \ne_47/ULTI1_33  ( .a(\ne_47/AEQB [33]), .b(\ne_47/LTV [33]), .out(
        \ne_47/LTV2 [33]) );
  nand2 \ne_47/ULTI2_33  ( .a(\ne_47/LTV1 [33]), .b(\ne_47/LTV2 [33]), .out(
        \ne_47/LTV [34]) );
  xor2 \ne_47/UEQI_34  ( .a(final_floor_elevator1[34]), .b(requested_floor[34]), .out(n2157) );
  nand2 \ne_47/UGTI0_34  ( .a(n2156), .b(final_floor_elevator1[34]), .out(
        \ne_47/GTV1 [34]) );
  nand2 \ne_47/UGTI1_34  ( .a(\ne_47/AEQB [34]), .b(\ne_47/GTV [34]), .out(
        \ne_47/GTV2 [34]) );
  nand2 \ne_47/UGTI2_34  ( .a(\ne_47/GTV1 [34]), .b(\ne_47/GTV2 [34]), .out(
        \ne_47/GTV [35]) );
  nand2 \ne_47/ULTI0_34  ( .a(n2155), .b(requested_floor[34]), .out(
        \ne_47/LTV1 [34]) );
  nand2 \ne_47/ULTI1_34  ( .a(\ne_47/AEQB [34]), .b(\ne_47/LTV [34]), .out(
        \ne_47/LTV2 [34]) );
  nand2 \ne_47/ULTI2_34  ( .a(\ne_47/LTV1 [34]), .b(\ne_47/LTV2 [34]), .out(
        \ne_47/LTV [35]) );
  xor2 \ne_47/UEQI_35  ( .a(final_floor_elevator1[35]), .b(requested_floor[35]), .out(n2154) );
  nand2 \ne_47/UGTI0_35  ( .a(n2153), .b(final_floor_elevator1[35]), .out(
        \ne_47/GTV1 [35]) );
  nand2 \ne_47/UGTI1_35  ( .a(\ne_47/AEQB [35]), .b(\ne_47/GTV [35]), .out(
        \ne_47/GTV2 [35]) );
  nand2 \ne_47/UGTI2_35  ( .a(\ne_47/GTV1 [35]), .b(\ne_47/GTV2 [35]), .out(
        \ne_47/GTV [36]) );
  nand2 \ne_47/ULTI0_35  ( .a(n2152), .b(requested_floor[35]), .out(
        \ne_47/LTV1 [35]) );
  nand2 \ne_47/ULTI1_35  ( .a(\ne_47/AEQB [35]), .b(\ne_47/LTV [35]), .out(
        \ne_47/LTV2 [35]) );
  nand2 \ne_47/ULTI2_35  ( .a(\ne_47/LTV1 [35]), .b(\ne_47/LTV2 [35]), .out(
        \ne_47/LTV [36]) );
  xor2 \ne_47/UEQI_36  ( .a(final_floor_elevator1[36]), .b(requested_floor[36]), .out(n2151) );
  nand2 \ne_47/UGTI0_36  ( .a(n2150), .b(final_floor_elevator1[36]), .out(
        \ne_47/GTV1 [36]) );
  nand2 \ne_47/UGTI1_36  ( .a(\ne_47/AEQB [36]), .b(\ne_47/GTV [36]), .out(
        \ne_47/GTV2 [36]) );
  nand2 \ne_47/UGTI2_36  ( .a(\ne_47/GTV1 [36]), .b(\ne_47/GTV2 [36]), .out(
        \ne_47/GTV [37]) );
  nand2 \ne_47/ULTI0_36  ( .a(n2149), .b(requested_floor[36]), .out(
        \ne_47/LTV1 [36]) );
  nand2 \ne_47/ULTI1_36  ( .a(\ne_47/AEQB [36]), .b(\ne_47/LTV [36]), .out(
        \ne_47/LTV2 [36]) );
  nand2 \ne_47/ULTI2_36  ( .a(\ne_47/LTV1 [36]), .b(\ne_47/LTV2 [36]), .out(
        \ne_47/LTV [37]) );
  xor2 \ne_47/UEQI_37  ( .a(final_floor_elevator1[37]), .b(requested_floor[37]), .out(n2148) );
  nand2 \ne_47/UGTI0_37  ( .a(n2147), .b(final_floor_elevator1[37]), .out(
        \ne_47/GTV1 [37]) );
  nand2 \ne_47/UGTI1_37  ( .a(\ne_47/AEQB [37]), .b(\ne_47/GTV [37]), .out(
        \ne_47/GTV2 [37]) );
  nand2 \ne_47/UGTI2_37  ( .a(\ne_47/GTV1 [37]), .b(\ne_47/GTV2 [37]), .out(
        \ne_47/GTV [38]) );
  nand2 \ne_47/ULTI0_37  ( .a(n2146), .b(requested_floor[37]), .out(
        \ne_47/LTV1 [37]) );
  nand2 \ne_47/ULTI1_37  ( .a(\ne_47/AEQB [37]), .b(\ne_47/LTV [37]), .out(
        \ne_47/LTV2 [37]) );
  nand2 \ne_47/ULTI2_37  ( .a(\ne_47/LTV1 [37]), .b(\ne_47/LTV2 [37]), .out(
        \ne_47/LTV [38]) );
  xor2 \ne_47/UEQI_38  ( .a(final_floor_elevator1[38]), .b(requested_floor[38]), .out(n2145) );
  nand2 \ne_47/UGTI0_38  ( .a(n2144), .b(final_floor_elevator1[38]), .out(
        \ne_47/GTV1 [38]) );
  nand2 \ne_47/UGTI1_38  ( .a(\ne_47/AEQB [38]), .b(\ne_47/GTV [38]), .out(
        \ne_47/GTV2 [38]) );
  nand2 \ne_47/UGTI2_38  ( .a(\ne_47/GTV1 [38]), .b(\ne_47/GTV2 [38]), .out(
        \ne_47/GTV [39]) );
  nand2 \ne_47/ULTI0_38  ( .a(n2143), .b(requested_floor[38]), .out(
        \ne_47/LTV1 [38]) );
  nand2 \ne_47/ULTI1_38  ( .a(\ne_47/AEQB [38]), .b(\ne_47/LTV [38]), .out(
        \ne_47/LTV2 [38]) );
  nand2 \ne_47/ULTI2_38  ( .a(\ne_47/LTV1 [38]), .b(\ne_47/LTV2 [38]), .out(
        \ne_47/LTV [39]) );
  xor2 \ne_47/UEQI_39  ( .a(final_floor_elevator1[39]), .b(requested_floor[39]), .out(n2142) );
  nand2 \ne_47/UGTI0_39  ( .a(n2141), .b(final_floor_elevator1[39]), .out(
        \ne_47/GTV1 [39]) );
  nand2 \ne_47/UGTI1_39  ( .a(\ne_47/AEQB [39]), .b(\ne_47/GTV [39]), .out(
        \ne_47/GTV2 [39]) );
  nand2 \ne_47/UGTI2_39  ( .a(\ne_47/GTV1 [39]), .b(\ne_47/GTV2 [39]), .out(
        \ne_47/GTV [40]) );
  nand2 \ne_47/ULTI0_39  ( .a(n2140), .b(requested_floor[39]), .out(
        \ne_47/LTV1 [39]) );
  nand2 \ne_47/ULTI1_39  ( .a(\ne_47/AEQB [39]), .b(\ne_47/LTV [39]), .out(
        \ne_47/LTV2 [39]) );
  nand2 \ne_47/ULTI2_39  ( .a(\ne_47/LTV1 [39]), .b(\ne_47/LTV2 [39]), .out(
        \ne_47/LTV [40]) );
  xor2 \ne_47/UEQI_40  ( .a(final_floor_elevator1[40]), .b(requested_floor[40]), .out(n2139) );
  nand2 \ne_47/UGTI0_40  ( .a(n2138), .b(final_floor_elevator1[40]), .out(
        \ne_47/GTV1 [40]) );
  nand2 \ne_47/UGTI1_40  ( .a(\ne_47/AEQB [40]), .b(\ne_47/GTV [40]), .out(
        \ne_47/GTV2 [40]) );
  nand2 \ne_47/UGTI2_40  ( .a(\ne_47/GTV1 [40]), .b(\ne_47/GTV2 [40]), .out(
        \ne_47/GTV [41]) );
  nand2 \ne_47/ULTI0_40  ( .a(n2137), .b(requested_floor[40]), .out(
        \ne_47/LTV1 [40]) );
  nand2 \ne_47/ULTI1_40  ( .a(\ne_47/AEQB [40]), .b(\ne_47/LTV [40]), .out(
        \ne_47/LTV2 [40]) );
  nand2 \ne_47/ULTI2_40  ( .a(\ne_47/LTV1 [40]), .b(\ne_47/LTV2 [40]), .out(
        \ne_47/LTV [41]) );
  xor2 \ne_47/UEQI_41  ( .a(final_floor_elevator1[41]), .b(requested_floor[41]), .out(n2136) );
  nand2 \ne_47/UGTI0_41  ( .a(n2135), .b(final_floor_elevator1[41]), .out(
        \ne_47/GTV1 [41]) );
  nand2 \ne_47/UGTI1_41  ( .a(\ne_47/AEQB [41]), .b(\ne_47/GTV [41]), .out(
        \ne_47/GTV2 [41]) );
  nand2 \ne_47/UGTI2_41  ( .a(\ne_47/GTV1 [41]), .b(\ne_47/GTV2 [41]), .out(
        \ne_47/GTV [42]) );
  nand2 \ne_47/ULTI0_41  ( .a(n2134), .b(requested_floor[41]), .out(
        \ne_47/LTV1 [41]) );
  nand2 \ne_47/ULTI1_41  ( .a(\ne_47/AEQB [41]), .b(\ne_47/LTV [41]), .out(
        \ne_47/LTV2 [41]) );
  nand2 \ne_47/ULTI2_41  ( .a(\ne_47/LTV1 [41]), .b(\ne_47/LTV2 [41]), .out(
        \ne_47/LTV [42]) );
  xor2 \ne_47/UEQI_42  ( .a(final_floor_elevator1[42]), .b(requested_floor[42]), .out(n2133) );
  nand2 \ne_47/UGTI0_42  ( .a(n2132), .b(final_floor_elevator1[42]), .out(
        \ne_47/GTV1 [42]) );
  nand2 \ne_47/UGTI1_42  ( .a(\ne_47/AEQB [42]), .b(\ne_47/GTV [42]), .out(
        \ne_47/GTV2 [42]) );
  nand2 \ne_47/UGTI2_42  ( .a(\ne_47/GTV1 [42]), .b(\ne_47/GTV2 [42]), .out(
        \ne_47/GTV [43]) );
  nand2 \ne_47/ULTI0_42  ( .a(n2131), .b(requested_floor[42]), .out(
        \ne_47/LTV1 [42]) );
  nand2 \ne_47/ULTI1_42  ( .a(\ne_47/AEQB [42]), .b(\ne_47/LTV [42]), .out(
        \ne_47/LTV2 [42]) );
  nand2 \ne_47/ULTI2_42  ( .a(\ne_47/LTV1 [42]), .b(\ne_47/LTV2 [42]), .out(
        \ne_47/LTV [43]) );
  xor2 \ne_47/UEQI_43  ( .a(final_floor_elevator1[43]), .b(requested_floor[43]), .out(n2130) );
  nand2 \ne_47/UGTI0_43  ( .a(n2129), .b(final_floor_elevator1[43]), .out(
        \ne_47/GTV1 [43]) );
  nand2 \ne_47/UGTI1_43  ( .a(\ne_47/AEQB [43]), .b(\ne_47/GTV [43]), .out(
        \ne_47/GTV2 [43]) );
  nand2 \ne_47/UGTI2_43  ( .a(\ne_47/GTV1 [43]), .b(\ne_47/GTV2 [43]), .out(
        \ne_47/GTV [44]) );
  nand2 \ne_47/ULTI0_43  ( .a(n2128), .b(requested_floor[43]), .out(
        \ne_47/LTV1 [43]) );
  nand2 \ne_47/ULTI1_43  ( .a(\ne_47/AEQB [43]), .b(\ne_47/LTV [43]), .out(
        \ne_47/LTV2 [43]) );
  nand2 \ne_47/ULTI2_43  ( .a(\ne_47/LTV1 [43]), .b(\ne_47/LTV2 [43]), .out(
        \ne_47/LTV [44]) );
  xor2 \ne_47/UEQI_44  ( .a(final_floor_elevator1[44]), .b(requested_floor[44]), .out(n2127) );
  nand2 \ne_47/UGTI0_44  ( .a(n2126), .b(final_floor_elevator1[44]), .out(
        \ne_47/GTV1 [44]) );
  nand2 \ne_47/UGTI1_44  ( .a(\ne_47/AEQB [44]), .b(\ne_47/GTV [44]), .out(
        \ne_47/GTV2 [44]) );
  nand2 \ne_47/UGTI2_44  ( .a(\ne_47/GTV1 [44]), .b(\ne_47/GTV2 [44]), .out(
        \ne_47/GTV [45]) );
  nand2 \ne_47/ULTI0_44  ( .a(n2125), .b(requested_floor[44]), .out(
        \ne_47/LTV1 [44]) );
  nand2 \ne_47/ULTI1_44  ( .a(\ne_47/AEQB [44]), .b(\ne_47/LTV [44]), .out(
        \ne_47/LTV2 [44]) );
  nand2 \ne_47/ULTI2_44  ( .a(\ne_47/LTV1 [44]), .b(\ne_47/LTV2 [44]), .out(
        \ne_47/LTV [45]) );
  xor2 \ne_47/UEQI_45  ( .a(final_floor_elevator1[45]), .b(requested_floor[45]), .out(n2124) );
  nand2 \ne_47/UGTI0_45  ( .a(n2123), .b(final_floor_elevator1[45]), .out(
        \ne_47/GTV1 [45]) );
  nand2 \ne_47/UGTI1_45  ( .a(\ne_47/AEQB [45]), .b(\ne_47/GTV [45]), .out(
        \ne_47/GTV2 [45]) );
  nand2 \ne_47/UGTI2_45  ( .a(\ne_47/GTV1 [45]), .b(\ne_47/GTV2 [45]), .out(
        \ne_47/GTV [46]) );
  nand2 \ne_47/ULTI0_45  ( .a(n2122), .b(requested_floor[45]), .out(
        \ne_47/LTV1 [45]) );
  nand2 \ne_47/ULTI1_45  ( .a(\ne_47/AEQB [45]), .b(\ne_47/LTV [45]), .out(
        \ne_47/LTV2 [45]) );
  nand2 \ne_47/ULTI2_45  ( .a(\ne_47/LTV1 [45]), .b(\ne_47/LTV2 [45]), .out(
        \ne_47/LTV [46]) );
  xor2 \ne_47/UEQI_46  ( .a(final_floor_elevator1[46]), .b(requested_floor[46]), .out(n2121) );
  nand2 \ne_47/UGTI0_46  ( .a(n2120), .b(final_floor_elevator1[46]), .out(
        \ne_47/GTV1 [46]) );
  nand2 \ne_47/UGTI1_46  ( .a(\ne_47/AEQB [46]), .b(\ne_47/GTV [46]), .out(
        \ne_47/GTV2 [46]) );
  nand2 \ne_47/UGTI2_46  ( .a(\ne_47/GTV1 [46]), .b(\ne_47/GTV2 [46]), .out(
        \ne_47/GTV [47]) );
  nand2 \ne_47/ULTI0_46  ( .a(n2119), .b(requested_floor[46]), .out(
        \ne_47/LTV1 [46]) );
  nand2 \ne_47/ULTI1_46  ( .a(\ne_47/AEQB [46]), .b(\ne_47/LTV [46]), .out(
        \ne_47/LTV2 [46]) );
  nand2 \ne_47/ULTI2_46  ( .a(\ne_47/LTV1 [46]), .b(\ne_47/LTV2 [46]), .out(
        \ne_47/LTV [47]) );
  xor2 \ne_47/UEQI_47  ( .a(final_floor_elevator1[47]), .b(requested_floor[47]), .out(n2118) );
  nand2 \ne_47/UGTI0_47  ( .a(n2117), .b(final_floor_elevator1[47]), .out(
        \ne_47/GTV1 [47]) );
  nand2 \ne_47/UGTI1_47  ( .a(\ne_47/AEQB [47]), .b(\ne_47/GTV [47]), .out(
        \ne_47/GTV2 [47]) );
  nand2 \ne_47/UGTI2_47  ( .a(\ne_47/GTV1 [47]), .b(\ne_47/GTV2 [47]), .out(
        \ne_47/GTV [48]) );
  nand2 \ne_47/ULTI0_47  ( .a(n2116), .b(requested_floor[47]), .out(
        \ne_47/LTV1 [47]) );
  nand2 \ne_47/ULTI1_47  ( .a(\ne_47/AEQB [47]), .b(\ne_47/LTV [47]), .out(
        \ne_47/LTV2 [47]) );
  nand2 \ne_47/ULTI2_47  ( .a(\ne_47/LTV1 [47]), .b(\ne_47/LTV2 [47]), .out(
        \ne_47/LTV [48]) );
  xor2 \ne_47/UEQI_48  ( .a(final_floor_elevator1[48]), .b(requested_floor[48]), .out(n2115) );
  nand2 \ne_47/UGTI0_48  ( .a(n2114), .b(final_floor_elevator1[48]), .out(
        \ne_47/GTV1 [48]) );
  nand2 \ne_47/UGTI1_48  ( .a(\ne_47/AEQB [48]), .b(\ne_47/GTV [48]), .out(
        \ne_47/GTV2 [48]) );
  nand2 \ne_47/UGTI2_48  ( .a(\ne_47/GTV1 [48]), .b(\ne_47/GTV2 [48]), .out(
        \ne_47/GTV [49]) );
  nand2 \ne_47/ULTI0_48  ( .a(n2113), .b(requested_floor[48]), .out(
        \ne_47/LTV1 [48]) );
  nand2 \ne_47/ULTI1_48  ( .a(\ne_47/AEQB [48]), .b(\ne_47/LTV [48]), .out(
        \ne_47/LTV2 [48]) );
  nand2 \ne_47/ULTI2_48  ( .a(\ne_47/LTV1 [48]), .b(\ne_47/LTV2 [48]), .out(
        \ne_47/LTV [49]) );
  xor2 \ne_47/UEQI_49  ( .a(final_floor_elevator1[49]), .b(requested_floor[49]), .out(n2112) );
  nand2 \ne_47/UGTI0_49  ( .a(n2111), .b(final_floor_elevator1[49]), .out(
        \ne_47/GTV1 [49]) );
  nand2 \ne_47/UGTI1_49  ( .a(\ne_47/AEQB [49]), .b(\ne_47/GTV [49]), .out(
        \ne_47/GTV2 [49]) );
  nand2 \ne_47/UGTI2_49  ( .a(\ne_47/GTV1 [49]), .b(\ne_47/GTV2 [49]), .out(
        \ne_47/GTV [50]) );
  nand2 \ne_47/ULTI0_49  ( .a(n2110), .b(requested_floor[49]), .out(
        \ne_47/LTV1 [49]) );
  nand2 \ne_47/ULTI1_49  ( .a(\ne_47/AEQB [49]), .b(\ne_47/LTV [49]), .out(
        \ne_47/LTV2 [49]) );
  nand2 \ne_47/ULTI2_49  ( .a(\ne_47/LTV1 [49]), .b(\ne_47/LTV2 [49]), .out(
        \ne_47/LTV [50]) );
  xor2 \ne_47/UEQI_50  ( .a(final_floor_elevator1[50]), .b(requested_floor[50]), .out(n2109) );
  nand2 \ne_47/UGTI0_50  ( .a(n2108), .b(final_floor_elevator1[50]), .out(
        \ne_47/GTV1 [50]) );
  nand2 \ne_47/UGTI1_50  ( .a(\ne_47/AEQB [50]), .b(\ne_47/GTV [50]), .out(
        \ne_47/GTV2 [50]) );
  nand2 \ne_47/UGTI2_50  ( .a(\ne_47/GTV1 [50]), .b(\ne_47/GTV2 [50]), .out(
        \ne_47/GTV [51]) );
  nand2 \ne_47/ULTI0_50  ( .a(n2107), .b(requested_floor[50]), .out(
        \ne_47/LTV1 [50]) );
  nand2 \ne_47/ULTI1_50  ( .a(\ne_47/AEQB [50]), .b(\ne_47/LTV [50]), .out(
        \ne_47/LTV2 [50]) );
  nand2 \ne_47/ULTI2_50  ( .a(\ne_47/LTV1 [50]), .b(\ne_47/LTV2 [50]), .out(
        \ne_47/LTV [51]) );
  xor2 \ne_47/UEQI_51  ( .a(final_floor_elevator1[51]), .b(requested_floor[51]), .out(n2106) );
  nand2 \ne_47/UGTI0_51  ( .a(n2105), .b(final_floor_elevator1[51]), .out(
        \ne_47/GTV1 [51]) );
  nand2 \ne_47/UGTI1_51  ( .a(\ne_47/AEQB [51]), .b(\ne_47/GTV [51]), .out(
        \ne_47/GTV2 [51]) );
  nand2 \ne_47/UGTI2_51  ( .a(\ne_47/GTV1 [51]), .b(\ne_47/GTV2 [51]), .out(
        \ne_47/GTV [52]) );
  nand2 \ne_47/ULTI0_51  ( .a(n2104), .b(requested_floor[51]), .out(
        \ne_47/LTV1 [51]) );
  nand2 \ne_47/ULTI1_51  ( .a(\ne_47/AEQB [51]), .b(\ne_47/LTV [51]), .out(
        \ne_47/LTV2 [51]) );
  nand2 \ne_47/ULTI2_51  ( .a(\ne_47/LTV1 [51]), .b(\ne_47/LTV2 [51]), .out(
        \ne_47/LTV [52]) );
  xor2 \ne_47/UEQI_52  ( .a(final_floor_elevator1[52]), .b(requested_floor[52]), .out(n2103) );
  nand2 \ne_47/UGTI0_52  ( .a(n2102), .b(final_floor_elevator1[52]), .out(
        \ne_47/GTV1 [52]) );
  nand2 \ne_47/UGTI1_52  ( .a(\ne_47/AEQB [52]), .b(\ne_47/GTV [52]), .out(
        \ne_47/GTV2 [52]) );
  nand2 \ne_47/UGTI2_52  ( .a(\ne_47/GTV1 [52]), .b(\ne_47/GTV2 [52]), .out(
        \ne_47/GTV [53]) );
  nand2 \ne_47/ULTI0_52  ( .a(n2101), .b(requested_floor[52]), .out(
        \ne_47/LTV1 [52]) );
  nand2 \ne_47/ULTI1_52  ( .a(\ne_47/AEQB [52]), .b(\ne_47/LTV [52]), .out(
        \ne_47/LTV2 [52]) );
  nand2 \ne_47/ULTI2_52  ( .a(\ne_47/LTV1 [52]), .b(\ne_47/LTV2 [52]), .out(
        \ne_47/LTV [53]) );
  xor2 \ne_47/UEQI_53  ( .a(final_floor_elevator1[53]), .b(requested_floor[53]), .out(n2100) );
  nand2 \ne_47/UGTI0_53  ( .a(n2099), .b(final_floor_elevator1[53]), .out(
        \ne_47/GTV1 [53]) );
  nand2 \ne_47/UGTI1_53  ( .a(\ne_47/AEQB [53]), .b(\ne_47/GTV [53]), .out(
        \ne_47/GTV2 [53]) );
  nand2 \ne_47/UGTI2_53  ( .a(\ne_47/GTV1 [53]), .b(\ne_47/GTV2 [53]), .out(
        \ne_47/GTV [54]) );
  nand2 \ne_47/ULTI0_53  ( .a(n2098), .b(requested_floor[53]), .out(
        \ne_47/LTV1 [53]) );
  nand2 \ne_47/ULTI1_53  ( .a(\ne_47/AEQB [53]), .b(\ne_47/LTV [53]), .out(
        \ne_47/LTV2 [53]) );
  nand2 \ne_47/ULTI2_53  ( .a(\ne_47/LTV1 [53]), .b(\ne_47/LTV2 [53]), .out(
        \ne_47/LTV [54]) );
  xor2 \ne_47/UEQI_54  ( .a(final_floor_elevator1[54]), .b(requested_floor[54]), .out(n2097) );
  nand2 \ne_47/UGTI0_54  ( .a(n2096), .b(final_floor_elevator1[54]), .out(
        \ne_47/GTV1 [54]) );
  nand2 \ne_47/UGTI1_54  ( .a(\ne_47/AEQB [54]), .b(\ne_47/GTV [54]), .out(
        \ne_47/GTV2 [54]) );
  nand2 \ne_47/UGTI2_54  ( .a(\ne_47/GTV1 [54]), .b(\ne_47/GTV2 [54]), .out(
        \ne_47/GTV [55]) );
  nand2 \ne_47/ULTI0_54  ( .a(n2095), .b(requested_floor[54]), .out(
        \ne_47/LTV1 [54]) );
  nand2 \ne_47/ULTI1_54  ( .a(\ne_47/AEQB [54]), .b(\ne_47/LTV [54]), .out(
        \ne_47/LTV2 [54]) );
  nand2 \ne_47/ULTI2_54  ( .a(\ne_47/LTV1 [54]), .b(\ne_47/LTV2 [54]), .out(
        \ne_47/LTV [55]) );
  xor2 \ne_47/UEQI_55  ( .a(final_floor_elevator1[55]), .b(requested_floor[55]), .out(n2094) );
  nand2 \ne_47/UGTI0_55  ( .a(n2093), .b(final_floor_elevator1[55]), .out(
        \ne_47/GTV1 [55]) );
  nand2 \ne_47/UGTI1_55  ( .a(\ne_47/AEQB [55]), .b(\ne_47/GTV [55]), .out(
        \ne_47/GTV2 [55]) );
  nand2 \ne_47/UGTI2_55  ( .a(\ne_47/GTV1 [55]), .b(\ne_47/GTV2 [55]), .out(
        \ne_47/GTV [56]) );
  nand2 \ne_47/ULTI0_55  ( .a(n2092), .b(requested_floor[55]), .out(
        \ne_47/LTV1 [55]) );
  nand2 \ne_47/ULTI1_55  ( .a(\ne_47/AEQB [55]), .b(\ne_47/LTV [55]), .out(
        \ne_47/LTV2 [55]) );
  nand2 \ne_47/ULTI2_55  ( .a(\ne_47/LTV1 [55]), .b(\ne_47/LTV2 [55]), .out(
        \ne_47/LTV [56]) );
  xor2 \ne_47/UEQI_56  ( .a(final_floor_elevator1[56]), .b(requested_floor[56]), .out(n2091) );
  nand2 \ne_47/UGTI0_56  ( .a(n2090), .b(final_floor_elevator1[56]), .out(
        \ne_47/GTV1 [56]) );
  nand2 \ne_47/UGTI1_56  ( .a(\ne_47/AEQB [56]), .b(\ne_47/GTV [56]), .out(
        \ne_47/GTV2 [56]) );
  nand2 \ne_47/UGTI2_56  ( .a(\ne_47/GTV1 [56]), .b(\ne_47/GTV2 [56]), .out(
        \ne_47/GTV [57]) );
  nand2 \ne_47/ULTI0_56  ( .a(n2089), .b(requested_floor[56]), .out(
        \ne_47/LTV1 [56]) );
  nand2 \ne_47/ULTI1_56  ( .a(\ne_47/AEQB [56]), .b(\ne_47/LTV [56]), .out(
        \ne_47/LTV2 [56]) );
  nand2 \ne_47/ULTI2_56  ( .a(\ne_47/LTV1 [56]), .b(\ne_47/LTV2 [56]), .out(
        \ne_47/LTV [57]) );
  xor2 \ne_47/UEQI_57  ( .a(final_floor_elevator1[57]), .b(requested_floor[57]), .out(n2088) );
  nand2 \ne_47/UGTI0_57  ( .a(n2087), .b(final_floor_elevator1[57]), .out(
        \ne_47/GTV1 [57]) );
  nand2 \ne_47/UGTI1_57  ( .a(\ne_47/AEQB [57]), .b(\ne_47/GTV [57]), .out(
        \ne_47/GTV2 [57]) );
  nand2 \ne_47/UGTI2_57  ( .a(\ne_47/GTV1 [57]), .b(\ne_47/GTV2 [57]), .out(
        \ne_47/GTV [58]) );
  nand2 \ne_47/ULTI0_57  ( .a(n2086), .b(requested_floor[57]), .out(
        \ne_47/LTV1 [57]) );
  nand2 \ne_47/ULTI1_57  ( .a(\ne_47/AEQB [57]), .b(\ne_47/LTV [57]), .out(
        \ne_47/LTV2 [57]) );
  nand2 \ne_47/ULTI2_57  ( .a(\ne_47/LTV1 [57]), .b(\ne_47/LTV2 [57]), .out(
        \ne_47/LTV [58]) );
  xor2 \ne_47/UEQI_58  ( .a(final_floor_elevator1[58]), .b(requested_floor[58]), .out(n2085) );
  nand2 \ne_47/UGTI0_58  ( .a(n2084), .b(final_floor_elevator1[58]), .out(
        \ne_47/GTV1 [58]) );
  nand2 \ne_47/UGTI1_58  ( .a(\ne_47/AEQB [58]), .b(\ne_47/GTV [58]), .out(
        \ne_47/GTV2 [58]) );
  nand2 \ne_47/UGTI2_58  ( .a(\ne_47/GTV1 [58]), .b(\ne_47/GTV2 [58]), .out(
        \ne_47/GTV [59]) );
  nand2 \ne_47/ULTI0_58  ( .a(n2083), .b(requested_floor[58]), .out(
        \ne_47/LTV1 [58]) );
  nand2 \ne_47/ULTI1_58  ( .a(\ne_47/AEQB [58]), .b(\ne_47/LTV [58]), .out(
        \ne_47/LTV2 [58]) );
  nand2 \ne_47/ULTI2_58  ( .a(\ne_47/LTV1 [58]), .b(\ne_47/LTV2 [58]), .out(
        \ne_47/LTV [59]) );
  xor2 \ne_47/UEQI_59  ( .a(final_floor_elevator1[59]), .b(requested_floor[59]), .out(n2082) );
  nand2 \ne_47/UGTI0_59  ( .a(n2081), .b(final_floor_elevator1[59]), .out(
        \ne_47/GTV1 [59]) );
  nand2 \ne_47/UGTI1_59  ( .a(\ne_47/AEQB [59]), .b(\ne_47/GTV [59]), .out(
        \ne_47/GTV2 [59]) );
  nand2 \ne_47/UGTI2_59  ( .a(\ne_47/GTV1 [59]), .b(\ne_47/GTV2 [59]), .out(
        \ne_47/GTV [60]) );
  nand2 \ne_47/ULTI0_59  ( .a(n2080), .b(requested_floor[59]), .out(
        \ne_47/LTV1 [59]) );
  nand2 \ne_47/ULTI1_59  ( .a(\ne_47/AEQB [59]), .b(\ne_47/LTV [59]), .out(
        \ne_47/LTV2 [59]) );
  nand2 \ne_47/ULTI2_59  ( .a(\ne_47/LTV1 [59]), .b(\ne_47/LTV2 [59]), .out(
        \ne_47/LTV [60]) );
  xor2 \ne_47/UEQI_60  ( .a(final_floor_elevator1[60]), .b(requested_floor[60]), .out(n2079) );
  nand2 \ne_47/UGTI0_60  ( .a(n2078), .b(final_floor_elevator1[60]), .out(
        \ne_47/GTV1 [60]) );
  nand2 \ne_47/UGTI1_60  ( .a(\ne_47/AEQB [60]), .b(\ne_47/GTV [60]), .out(
        \ne_47/GTV2 [60]) );
  nand2 \ne_47/UGTI2_60  ( .a(\ne_47/GTV1 [60]), .b(\ne_47/GTV2 [60]), .out(
        \ne_47/GTV [61]) );
  nand2 \ne_47/ULTI0_60  ( .a(n2077), .b(requested_floor[60]), .out(
        \ne_47/LTV1 [60]) );
  nand2 \ne_47/ULTI1_60  ( .a(\ne_47/AEQB [60]), .b(\ne_47/LTV [60]), .out(
        \ne_47/LTV2 [60]) );
  nand2 \ne_47/ULTI2_60  ( .a(\ne_47/LTV1 [60]), .b(\ne_47/LTV2 [60]), .out(
        \ne_47/LTV [61]) );
  xor2 \ne_47/UEQI_61  ( .a(final_floor_elevator1[61]), .b(requested_floor[61]), .out(n2076) );
  nand2 \ne_47/UGTI0_61  ( .a(n2075), .b(final_floor_elevator1[61]), .out(
        \ne_47/GTV1 [61]) );
  nand2 \ne_47/UGTI1_61  ( .a(\ne_47/AEQB [61]), .b(\ne_47/GTV [61]), .out(
        \ne_47/GTV2 [61]) );
  nand2 \ne_47/UGTI2_61  ( .a(\ne_47/GTV1 [61]), .b(\ne_47/GTV2 [61]), .out(
        \ne_47/GTV [62]) );
  nand2 \ne_47/ULTI0_61  ( .a(n2074), .b(requested_floor[61]), .out(
        \ne_47/LTV1 [61]) );
  nand2 \ne_47/ULTI1_61  ( .a(\ne_47/AEQB [61]), .b(\ne_47/LTV [61]), .out(
        \ne_47/LTV2 [61]) );
  nand2 \ne_47/ULTI2_61  ( .a(\ne_47/LTV1 [61]), .b(\ne_47/LTV2 [61]), .out(
        \ne_47/LTV [62]) );
  xor2 \ne_47/UEQI_62  ( .a(final_floor_elevator1[62]), .b(requested_floor[62]), .out(n2073) );
  nand2 \ne_47/UGTI0_62  ( .a(n2072), .b(final_floor_elevator1[62]), .out(
        \ne_47/GTV1 [62]) );
  nand2 \ne_47/UGTI1_62  ( .a(\ne_47/AEQB [62]), .b(\ne_47/GTV [62]), .out(
        \ne_47/GTV2 [62]) );
  nand2 \ne_47/UGTI2_62  ( .a(\ne_47/GTV1 [62]), .b(\ne_47/GTV2 [62]), .out(
        \ne_47/GTV [63]) );
  nand2 \ne_47/ULTI0_62  ( .a(n2071), .b(requested_floor[62]), .out(
        \ne_47/LTV1 [62]) );
  nand2 \ne_47/ULTI1_62  ( .a(\ne_47/AEQB [62]), .b(\ne_47/LTV [62]), .out(
        \ne_47/LTV2 [62]) );
  nand2 \ne_47/ULTI2_62  ( .a(\ne_47/LTV1 [62]), .b(\ne_47/LTV2 [62]), .out(
        \ne_47/LTV [63]) );
  nor2 \eq_42_3/UEQ  ( .a(\eq_42_3/GT ), .b(\eq_42_3/LT ), .out(N13) );
  nand2 \eq_42_3/UNGT0  ( .a(current_floor_output_elevator1[0]), .b(n2070), 
        .out(n2069) );
  nand2 \eq_42_3/UNLT0  ( .a(destination_floor_elevator1[0]), .b(n2068), .out(
        n2067) );
  xor2 \eq_42_3/UEQI  ( .a(\eq_42_3/SA ), .b(\eq_42_3/SB ), .out(n2066) );
  nand2 \eq_42_3/UGTI0  ( .a(n2065), .b(\eq_42_3/SA ), .out(\eq_42_3/GTV1 [63]) );
  nand2 \eq_42_3/UGTI1  ( .a(\eq_42_3/AEQB [63]), .b(\eq_42_3/GTV [63]), .out(
        \eq_42_3/GTV2 [63]) );
  nand2 \eq_42_3/UGTI2  ( .a(\eq_42_3/GTV1 [63]), .b(\eq_42_3/GTV2 [63]), 
        .out(\eq_42_3/GT ) );
  nand2 \eq_42_3/ULTI0  ( .a(n2064), .b(\eq_42_3/SB ), .out(\eq_42_3/LTV1 [63]) );
  nand2 \eq_42_3/ULTI1  ( .a(\eq_42_3/AEQB [63]), .b(\eq_42_3/LTV [63]), .out(
        \eq_42_3/LTV2 [63]) );
  nand2 \eq_42_3/ULTI2  ( .a(\eq_42_3/LTV1 [63]), .b(\eq_42_3/LTV2 [63]), 
        .out(\eq_42_3/LT ) );
  xor2 \eq_42_3/UEQI_1  ( .a(current_floor_output_elevator1[1]), .b(
        destination_floor_elevator1[1]), .out(n2063) );
  nand2 \eq_42_3/UGTI0_1  ( .a(n2062), .b(current_floor_output_elevator1[1]), 
        .out(\eq_42_3/GTV1 [1]) );
  nand2 \eq_42_3/UGTI1_1  ( .a(\eq_42_3/AEQB [1]), .b(\eq_42_3/GTV [1]), .out(
        \eq_42_3/GTV2 [1]) );
  nand2 \eq_42_3/UGTI2_1  ( .a(\eq_42_3/GTV1 [1]), .b(\eq_42_3/GTV2 [1]), 
        .out(\eq_42_3/GTV [2]) );
  nand2 \eq_42_3/ULTI0_1  ( .a(n2061), .b(destination_floor_elevator1[1]), 
        .out(\eq_42_3/LTV1 [1]) );
  nand2 \eq_42_3/ULTI1_1  ( .a(\eq_42_3/AEQB [1]), .b(\eq_42_3/LTV [1]), .out(
        \eq_42_3/LTV2 [1]) );
  nand2 \eq_42_3/ULTI2_1  ( .a(\eq_42_3/LTV1 [1]), .b(\eq_42_3/LTV2 [1]), 
        .out(\eq_42_3/LTV [2]) );
  xor2 \eq_42_3/UEQI_2  ( .a(current_floor_output_elevator1[2]), .b(
        destination_floor_elevator1[2]), .out(n2060) );
  nand2 \eq_42_3/UGTI0_2  ( .a(n2059), .b(current_floor_output_elevator1[2]), 
        .out(\eq_42_3/GTV1 [2]) );
  nand2 \eq_42_3/UGTI1_2  ( .a(\eq_42_3/AEQB [2]), .b(\eq_42_3/GTV [2]), .out(
        \eq_42_3/GTV2 [2]) );
  nand2 \eq_42_3/UGTI2_2  ( .a(\eq_42_3/GTV1 [2]), .b(\eq_42_3/GTV2 [2]), 
        .out(\eq_42_3/GTV [3]) );
  nand2 \eq_42_3/ULTI0_2  ( .a(n2058), .b(destination_floor_elevator1[2]), 
        .out(\eq_42_3/LTV1 [2]) );
  nand2 \eq_42_3/ULTI1_2  ( .a(\eq_42_3/AEQB [2]), .b(\eq_42_3/LTV [2]), .out(
        \eq_42_3/LTV2 [2]) );
  nand2 \eq_42_3/ULTI2_2  ( .a(\eq_42_3/LTV1 [2]), .b(\eq_42_3/LTV2 [2]), 
        .out(\eq_42_3/LTV [3]) );
  xor2 \eq_42_3/UEQI_3  ( .a(current_floor_output_elevator1[3]), .b(
        destination_floor_elevator1[3]), .out(n2057) );
  nand2 \eq_42_3/UGTI0_3  ( .a(n2056), .b(current_floor_output_elevator1[3]), 
        .out(\eq_42_3/GTV1 [3]) );
  nand2 \eq_42_3/UGTI1_3  ( .a(\eq_42_3/AEQB [3]), .b(\eq_42_3/GTV [3]), .out(
        \eq_42_3/GTV2 [3]) );
  nand2 \eq_42_3/UGTI2_3  ( .a(\eq_42_3/GTV1 [3]), .b(\eq_42_3/GTV2 [3]), 
        .out(\eq_42_3/GTV [4]) );
  nand2 \eq_42_3/ULTI0_3  ( .a(n2055), .b(destination_floor_elevator1[3]), 
        .out(\eq_42_3/LTV1 [3]) );
  nand2 \eq_42_3/ULTI1_3  ( .a(\eq_42_3/AEQB [3]), .b(\eq_42_3/LTV [3]), .out(
        \eq_42_3/LTV2 [3]) );
  nand2 \eq_42_3/ULTI2_3  ( .a(\eq_42_3/LTV1 [3]), .b(\eq_42_3/LTV2 [3]), 
        .out(\eq_42_3/LTV [4]) );
  xor2 \eq_42_3/UEQI_4  ( .a(current_floor_output_elevator1[4]), .b(
        destination_floor_elevator1[4]), .out(n2054) );
  nand2 \eq_42_3/UGTI0_4  ( .a(n2053), .b(current_floor_output_elevator1[4]), 
        .out(\eq_42_3/GTV1 [4]) );
  nand2 \eq_42_3/UGTI1_4  ( .a(\eq_42_3/AEQB [4]), .b(\eq_42_3/GTV [4]), .out(
        \eq_42_3/GTV2 [4]) );
  nand2 \eq_42_3/UGTI2_4  ( .a(\eq_42_3/GTV1 [4]), .b(\eq_42_3/GTV2 [4]), 
        .out(\eq_42_3/GTV [5]) );
  nand2 \eq_42_3/ULTI0_4  ( .a(n2052), .b(destination_floor_elevator1[4]), 
        .out(\eq_42_3/LTV1 [4]) );
  nand2 \eq_42_3/ULTI1_4  ( .a(\eq_42_3/AEQB [4]), .b(\eq_42_3/LTV [4]), .out(
        \eq_42_3/LTV2 [4]) );
  nand2 \eq_42_3/ULTI2_4  ( .a(\eq_42_3/LTV1 [4]), .b(\eq_42_3/LTV2 [4]), 
        .out(\eq_42_3/LTV [5]) );
  xor2 \eq_42_3/UEQI_5  ( .a(current_floor_output_elevator1[5]), .b(
        destination_floor_elevator1[5]), .out(n2051) );
  nand2 \eq_42_3/UGTI0_5  ( .a(n2050), .b(current_floor_output_elevator1[5]), 
        .out(\eq_42_3/GTV1 [5]) );
  nand2 \eq_42_3/UGTI1_5  ( .a(\eq_42_3/AEQB [5]), .b(\eq_42_3/GTV [5]), .out(
        \eq_42_3/GTV2 [5]) );
  nand2 \eq_42_3/UGTI2_5  ( .a(\eq_42_3/GTV1 [5]), .b(\eq_42_3/GTV2 [5]), 
        .out(\eq_42_3/GTV [6]) );
  nand2 \eq_42_3/ULTI0_5  ( .a(n2049), .b(destination_floor_elevator1[5]), 
        .out(\eq_42_3/LTV1 [5]) );
  nand2 \eq_42_3/ULTI1_5  ( .a(\eq_42_3/AEQB [5]), .b(\eq_42_3/LTV [5]), .out(
        \eq_42_3/LTV2 [5]) );
  nand2 \eq_42_3/ULTI2_5  ( .a(\eq_42_3/LTV1 [5]), .b(\eq_42_3/LTV2 [5]), 
        .out(\eq_42_3/LTV [6]) );
  xor2 \eq_42_3/UEQI_6  ( .a(current_floor_output_elevator1[6]), .b(
        destination_floor_elevator1[6]), .out(n2048) );
  nand2 \eq_42_3/UGTI0_6  ( .a(n2047), .b(current_floor_output_elevator1[6]), 
        .out(\eq_42_3/GTV1 [6]) );
  nand2 \eq_42_3/UGTI1_6  ( .a(\eq_42_3/AEQB [6]), .b(\eq_42_3/GTV [6]), .out(
        \eq_42_3/GTV2 [6]) );
  nand2 \eq_42_3/UGTI2_6  ( .a(\eq_42_3/GTV1 [6]), .b(\eq_42_3/GTV2 [6]), 
        .out(\eq_42_3/GTV [7]) );
  nand2 \eq_42_3/ULTI0_6  ( .a(n2046), .b(destination_floor_elevator1[6]), 
        .out(\eq_42_3/LTV1 [6]) );
  nand2 \eq_42_3/ULTI1_6  ( .a(\eq_42_3/AEQB [6]), .b(\eq_42_3/LTV [6]), .out(
        \eq_42_3/LTV2 [6]) );
  nand2 \eq_42_3/ULTI2_6  ( .a(\eq_42_3/LTV1 [6]), .b(\eq_42_3/LTV2 [6]), 
        .out(\eq_42_3/LTV [7]) );
  xor2 \eq_42_3/UEQI_7  ( .a(current_floor_output_elevator1[7]), .b(
        destination_floor_elevator1[7]), .out(n2045) );
  nand2 \eq_42_3/UGTI0_7  ( .a(n2044), .b(current_floor_output_elevator1[7]), 
        .out(\eq_42_3/GTV1 [7]) );
  nand2 \eq_42_3/UGTI1_7  ( .a(\eq_42_3/AEQB [7]), .b(\eq_42_3/GTV [7]), .out(
        \eq_42_3/GTV2 [7]) );
  nand2 \eq_42_3/UGTI2_7  ( .a(\eq_42_3/GTV1 [7]), .b(\eq_42_3/GTV2 [7]), 
        .out(\eq_42_3/GTV [8]) );
  nand2 \eq_42_3/ULTI0_7  ( .a(n2043), .b(destination_floor_elevator1[7]), 
        .out(\eq_42_3/LTV1 [7]) );
  nand2 \eq_42_3/ULTI1_7  ( .a(\eq_42_3/AEQB [7]), .b(\eq_42_3/LTV [7]), .out(
        \eq_42_3/LTV2 [7]) );
  nand2 \eq_42_3/ULTI2_7  ( .a(\eq_42_3/LTV1 [7]), .b(\eq_42_3/LTV2 [7]), 
        .out(\eq_42_3/LTV [8]) );
  xor2 \eq_42_3/UEQI_8  ( .a(current_floor_output_elevator1[8]), .b(
        destination_floor_elevator1[8]), .out(n2042) );
  nand2 \eq_42_3/UGTI0_8  ( .a(n2041), .b(current_floor_output_elevator1[8]), 
        .out(\eq_42_3/GTV1 [8]) );
  nand2 \eq_42_3/UGTI1_8  ( .a(\eq_42_3/AEQB [8]), .b(\eq_42_3/GTV [8]), .out(
        \eq_42_3/GTV2 [8]) );
  nand2 \eq_42_3/UGTI2_8  ( .a(\eq_42_3/GTV1 [8]), .b(\eq_42_3/GTV2 [8]), 
        .out(\eq_42_3/GTV [9]) );
  nand2 \eq_42_3/ULTI0_8  ( .a(n2040), .b(destination_floor_elevator1[8]), 
        .out(\eq_42_3/LTV1 [8]) );
  nand2 \eq_42_3/ULTI1_8  ( .a(\eq_42_3/AEQB [8]), .b(\eq_42_3/LTV [8]), .out(
        \eq_42_3/LTV2 [8]) );
  nand2 \eq_42_3/ULTI2_8  ( .a(\eq_42_3/LTV1 [8]), .b(\eq_42_3/LTV2 [8]), 
        .out(\eq_42_3/LTV [9]) );
  xor2 \eq_42_3/UEQI_9  ( .a(current_floor_output_elevator1[9]), .b(
        destination_floor_elevator1[9]), .out(n2039) );
  nand2 \eq_42_3/UGTI0_9  ( .a(n2038), .b(current_floor_output_elevator1[9]), 
        .out(\eq_42_3/GTV1 [9]) );
  nand2 \eq_42_3/UGTI1_9  ( .a(\eq_42_3/AEQB [9]), .b(\eq_42_3/GTV [9]), .out(
        \eq_42_3/GTV2 [9]) );
  nand2 \eq_42_3/UGTI2_9  ( .a(\eq_42_3/GTV1 [9]), .b(\eq_42_3/GTV2 [9]), 
        .out(\eq_42_3/GTV [10]) );
  nand2 \eq_42_3/ULTI0_9  ( .a(n2037), .b(destination_floor_elevator1[9]), 
        .out(\eq_42_3/LTV1 [9]) );
  nand2 \eq_42_3/ULTI1_9  ( .a(\eq_42_3/AEQB [9]), .b(\eq_42_3/LTV [9]), .out(
        \eq_42_3/LTV2 [9]) );
  nand2 \eq_42_3/ULTI2_9  ( .a(\eq_42_3/LTV1 [9]), .b(\eq_42_3/LTV2 [9]), 
        .out(\eq_42_3/LTV [10]) );
  xor2 \eq_42_3/UEQI_10  ( .a(current_floor_output_elevator1[10]), .b(
        destination_floor_elevator1[10]), .out(n2036) );
  nand2 \eq_42_3/UGTI0_10  ( .a(n2035), .b(current_floor_output_elevator1[10]), 
        .out(\eq_42_3/GTV1 [10]) );
  nand2 \eq_42_3/UGTI1_10  ( .a(\eq_42_3/AEQB [10]), .b(\eq_42_3/GTV [10]), 
        .out(\eq_42_3/GTV2 [10]) );
  nand2 \eq_42_3/UGTI2_10  ( .a(\eq_42_3/GTV1 [10]), .b(\eq_42_3/GTV2 [10]), 
        .out(\eq_42_3/GTV [11]) );
  nand2 \eq_42_3/ULTI0_10  ( .a(n2034), .b(destination_floor_elevator1[10]), 
        .out(\eq_42_3/LTV1 [10]) );
  nand2 \eq_42_3/ULTI1_10  ( .a(\eq_42_3/AEQB [10]), .b(\eq_42_3/LTV [10]), 
        .out(\eq_42_3/LTV2 [10]) );
  nand2 \eq_42_3/ULTI2_10  ( .a(\eq_42_3/LTV1 [10]), .b(\eq_42_3/LTV2 [10]), 
        .out(\eq_42_3/LTV [11]) );
  xor2 \eq_42_3/UEQI_11  ( .a(current_floor_output_elevator1[11]), .b(
        destination_floor_elevator1[11]), .out(n2033) );
  nand2 \eq_42_3/UGTI0_11  ( .a(n2032), .b(current_floor_output_elevator1[11]), 
        .out(\eq_42_3/GTV1 [11]) );
  nand2 \eq_42_3/UGTI1_11  ( .a(\eq_42_3/AEQB [11]), .b(\eq_42_3/GTV [11]), 
        .out(\eq_42_3/GTV2 [11]) );
  nand2 \eq_42_3/UGTI2_11  ( .a(\eq_42_3/GTV1 [11]), .b(\eq_42_3/GTV2 [11]), 
        .out(\eq_42_3/GTV [12]) );
  nand2 \eq_42_3/ULTI0_11  ( .a(n2031), .b(destination_floor_elevator1[11]), 
        .out(\eq_42_3/LTV1 [11]) );
  nand2 \eq_42_3/ULTI1_11  ( .a(\eq_42_3/AEQB [11]), .b(\eq_42_3/LTV [11]), 
        .out(\eq_42_3/LTV2 [11]) );
  nand2 \eq_42_3/ULTI2_11  ( .a(\eq_42_3/LTV1 [11]), .b(\eq_42_3/LTV2 [11]), 
        .out(\eq_42_3/LTV [12]) );
  xor2 \eq_42_3/UEQI_12  ( .a(current_floor_output_elevator1[12]), .b(
        destination_floor_elevator1[12]), .out(n2030) );
  nand2 \eq_42_3/UGTI0_12  ( .a(n2029), .b(current_floor_output_elevator1[12]), 
        .out(\eq_42_3/GTV1 [12]) );
  nand2 \eq_42_3/UGTI1_12  ( .a(\eq_42_3/AEQB [12]), .b(\eq_42_3/GTV [12]), 
        .out(\eq_42_3/GTV2 [12]) );
  nand2 \eq_42_3/UGTI2_12  ( .a(\eq_42_3/GTV1 [12]), .b(\eq_42_3/GTV2 [12]), 
        .out(\eq_42_3/GTV [13]) );
  nand2 \eq_42_3/ULTI0_12  ( .a(n2028), .b(destination_floor_elevator1[12]), 
        .out(\eq_42_3/LTV1 [12]) );
  nand2 \eq_42_3/ULTI1_12  ( .a(\eq_42_3/AEQB [12]), .b(\eq_42_3/LTV [12]), 
        .out(\eq_42_3/LTV2 [12]) );
  nand2 \eq_42_3/ULTI2_12  ( .a(\eq_42_3/LTV1 [12]), .b(\eq_42_3/LTV2 [12]), 
        .out(\eq_42_3/LTV [13]) );
  xor2 \eq_42_3/UEQI_13  ( .a(current_floor_output_elevator1[13]), .b(
        destination_floor_elevator1[13]), .out(n2027) );
  nand2 \eq_42_3/UGTI0_13  ( .a(n2026), .b(current_floor_output_elevator1[13]), 
        .out(\eq_42_3/GTV1 [13]) );
  nand2 \eq_42_3/UGTI1_13  ( .a(\eq_42_3/AEQB [13]), .b(\eq_42_3/GTV [13]), 
        .out(\eq_42_3/GTV2 [13]) );
  nand2 \eq_42_3/UGTI2_13  ( .a(\eq_42_3/GTV1 [13]), .b(\eq_42_3/GTV2 [13]), 
        .out(\eq_42_3/GTV [14]) );
  nand2 \eq_42_3/ULTI0_13  ( .a(n2025), .b(destination_floor_elevator1[13]), 
        .out(\eq_42_3/LTV1 [13]) );
  nand2 \eq_42_3/ULTI1_13  ( .a(\eq_42_3/AEQB [13]), .b(\eq_42_3/LTV [13]), 
        .out(\eq_42_3/LTV2 [13]) );
  nand2 \eq_42_3/ULTI2_13  ( .a(\eq_42_3/LTV1 [13]), .b(\eq_42_3/LTV2 [13]), 
        .out(\eq_42_3/LTV [14]) );
  xor2 \eq_42_3/UEQI_14  ( .a(current_floor_output_elevator1[14]), .b(
        destination_floor_elevator1[14]), .out(n2024) );
  nand2 \eq_42_3/UGTI0_14  ( .a(n2023), .b(current_floor_output_elevator1[14]), 
        .out(\eq_42_3/GTV1 [14]) );
  nand2 \eq_42_3/UGTI1_14  ( .a(\eq_42_3/AEQB [14]), .b(\eq_42_3/GTV [14]), 
        .out(\eq_42_3/GTV2 [14]) );
  nand2 \eq_42_3/UGTI2_14  ( .a(\eq_42_3/GTV1 [14]), .b(\eq_42_3/GTV2 [14]), 
        .out(\eq_42_3/GTV [15]) );
  nand2 \eq_42_3/ULTI0_14  ( .a(n2022), .b(destination_floor_elevator1[14]), 
        .out(\eq_42_3/LTV1 [14]) );
  nand2 \eq_42_3/ULTI1_14  ( .a(\eq_42_3/AEQB [14]), .b(\eq_42_3/LTV [14]), 
        .out(\eq_42_3/LTV2 [14]) );
  nand2 \eq_42_3/ULTI2_14  ( .a(\eq_42_3/LTV1 [14]), .b(\eq_42_3/LTV2 [14]), 
        .out(\eq_42_3/LTV [15]) );
  xor2 \eq_42_3/UEQI_15  ( .a(current_floor_output_elevator1[15]), .b(
        destination_floor_elevator1[15]), .out(n2021) );
  nand2 \eq_42_3/UGTI0_15  ( .a(n2020), .b(current_floor_output_elevator1[15]), 
        .out(\eq_42_3/GTV1 [15]) );
  nand2 \eq_42_3/UGTI1_15  ( .a(\eq_42_3/AEQB [15]), .b(\eq_42_3/GTV [15]), 
        .out(\eq_42_3/GTV2 [15]) );
  nand2 \eq_42_3/UGTI2_15  ( .a(\eq_42_3/GTV1 [15]), .b(\eq_42_3/GTV2 [15]), 
        .out(\eq_42_3/GTV [16]) );
  nand2 \eq_42_3/ULTI0_15  ( .a(n2019), .b(destination_floor_elevator1[15]), 
        .out(\eq_42_3/LTV1 [15]) );
  nand2 \eq_42_3/ULTI1_15  ( .a(\eq_42_3/AEQB [15]), .b(\eq_42_3/LTV [15]), 
        .out(\eq_42_3/LTV2 [15]) );
  nand2 \eq_42_3/ULTI2_15  ( .a(\eq_42_3/LTV1 [15]), .b(\eq_42_3/LTV2 [15]), 
        .out(\eq_42_3/LTV [16]) );
  xor2 \eq_42_3/UEQI_16  ( .a(current_floor_output_elevator1[16]), .b(
        destination_floor_elevator1[16]), .out(n2018) );
  nand2 \eq_42_3/UGTI0_16  ( .a(n2017), .b(current_floor_output_elevator1[16]), 
        .out(\eq_42_3/GTV1 [16]) );
  nand2 \eq_42_3/UGTI1_16  ( .a(\eq_42_3/AEQB [16]), .b(\eq_42_3/GTV [16]), 
        .out(\eq_42_3/GTV2 [16]) );
  nand2 \eq_42_3/UGTI2_16  ( .a(\eq_42_3/GTV1 [16]), .b(\eq_42_3/GTV2 [16]), 
        .out(\eq_42_3/GTV [17]) );
  nand2 \eq_42_3/ULTI0_16  ( .a(n2016), .b(destination_floor_elevator1[16]), 
        .out(\eq_42_3/LTV1 [16]) );
  nand2 \eq_42_3/ULTI1_16  ( .a(\eq_42_3/AEQB [16]), .b(\eq_42_3/LTV [16]), 
        .out(\eq_42_3/LTV2 [16]) );
  nand2 \eq_42_3/ULTI2_16  ( .a(\eq_42_3/LTV1 [16]), .b(\eq_42_3/LTV2 [16]), 
        .out(\eq_42_3/LTV [17]) );
  xor2 \eq_42_3/UEQI_17  ( .a(current_floor_output_elevator1[17]), .b(
        destination_floor_elevator1[17]), .out(n2015) );
  nand2 \eq_42_3/UGTI0_17  ( .a(n2014), .b(current_floor_output_elevator1[17]), 
        .out(\eq_42_3/GTV1 [17]) );
  nand2 \eq_42_3/UGTI1_17  ( .a(\eq_42_3/AEQB [17]), .b(\eq_42_3/GTV [17]), 
        .out(\eq_42_3/GTV2 [17]) );
  nand2 \eq_42_3/UGTI2_17  ( .a(\eq_42_3/GTV1 [17]), .b(\eq_42_3/GTV2 [17]), 
        .out(\eq_42_3/GTV [18]) );
  nand2 \eq_42_3/ULTI0_17  ( .a(n2013), .b(destination_floor_elevator1[17]), 
        .out(\eq_42_3/LTV1 [17]) );
  nand2 \eq_42_3/ULTI1_17  ( .a(\eq_42_3/AEQB [17]), .b(\eq_42_3/LTV [17]), 
        .out(\eq_42_3/LTV2 [17]) );
  nand2 \eq_42_3/ULTI2_17  ( .a(\eq_42_3/LTV1 [17]), .b(\eq_42_3/LTV2 [17]), 
        .out(\eq_42_3/LTV [18]) );
  xor2 \eq_42_3/UEQI_18  ( .a(current_floor_output_elevator1[18]), .b(
        destination_floor_elevator1[18]), .out(n2012) );
  nand2 \eq_42_3/UGTI0_18  ( .a(n2011), .b(current_floor_output_elevator1[18]), 
        .out(\eq_42_3/GTV1 [18]) );
  nand2 \eq_42_3/UGTI1_18  ( .a(\eq_42_3/AEQB [18]), .b(\eq_42_3/GTV [18]), 
        .out(\eq_42_3/GTV2 [18]) );
  nand2 \eq_42_3/UGTI2_18  ( .a(\eq_42_3/GTV1 [18]), .b(\eq_42_3/GTV2 [18]), 
        .out(\eq_42_3/GTV [19]) );
  nand2 \eq_42_3/ULTI0_18  ( .a(n2010), .b(destination_floor_elevator1[18]), 
        .out(\eq_42_3/LTV1 [18]) );
  nand2 \eq_42_3/ULTI1_18  ( .a(\eq_42_3/AEQB [18]), .b(\eq_42_3/LTV [18]), 
        .out(\eq_42_3/LTV2 [18]) );
  nand2 \eq_42_3/ULTI2_18  ( .a(\eq_42_3/LTV1 [18]), .b(\eq_42_3/LTV2 [18]), 
        .out(\eq_42_3/LTV [19]) );
  xor2 \eq_42_3/UEQI_19  ( .a(current_floor_output_elevator1[19]), .b(
        destination_floor_elevator1[19]), .out(n2009) );
  nand2 \eq_42_3/UGTI0_19  ( .a(n2008), .b(current_floor_output_elevator1[19]), 
        .out(\eq_42_3/GTV1 [19]) );
  nand2 \eq_42_3/UGTI1_19  ( .a(\eq_42_3/AEQB [19]), .b(\eq_42_3/GTV [19]), 
        .out(\eq_42_3/GTV2 [19]) );
  nand2 \eq_42_3/UGTI2_19  ( .a(\eq_42_3/GTV1 [19]), .b(\eq_42_3/GTV2 [19]), 
        .out(\eq_42_3/GTV [20]) );
  nand2 \eq_42_3/ULTI0_19  ( .a(n2007), .b(destination_floor_elevator1[19]), 
        .out(\eq_42_3/LTV1 [19]) );
  nand2 \eq_42_3/ULTI1_19  ( .a(\eq_42_3/AEQB [19]), .b(\eq_42_3/LTV [19]), 
        .out(\eq_42_3/LTV2 [19]) );
  nand2 \eq_42_3/ULTI2_19  ( .a(\eq_42_3/LTV1 [19]), .b(\eq_42_3/LTV2 [19]), 
        .out(\eq_42_3/LTV [20]) );
  xor2 \eq_42_3/UEQI_20  ( .a(current_floor_output_elevator1[20]), .b(
        destination_floor_elevator1[20]), .out(n2006) );
  nand2 \eq_42_3/UGTI0_20  ( .a(n2005), .b(current_floor_output_elevator1[20]), 
        .out(\eq_42_3/GTV1 [20]) );
  nand2 \eq_42_3/UGTI1_20  ( .a(\eq_42_3/AEQB [20]), .b(\eq_42_3/GTV [20]), 
        .out(\eq_42_3/GTV2 [20]) );
  nand2 \eq_42_3/UGTI2_20  ( .a(\eq_42_3/GTV1 [20]), .b(\eq_42_3/GTV2 [20]), 
        .out(\eq_42_3/GTV [21]) );
  nand2 \eq_42_3/ULTI0_20  ( .a(n2004), .b(destination_floor_elevator1[20]), 
        .out(\eq_42_3/LTV1 [20]) );
  nand2 \eq_42_3/ULTI1_20  ( .a(\eq_42_3/AEQB [20]), .b(\eq_42_3/LTV [20]), 
        .out(\eq_42_3/LTV2 [20]) );
  nand2 \eq_42_3/ULTI2_20  ( .a(\eq_42_3/LTV1 [20]), .b(\eq_42_3/LTV2 [20]), 
        .out(\eq_42_3/LTV [21]) );
  xor2 \eq_42_3/UEQI_21  ( .a(current_floor_output_elevator1[21]), .b(
        destination_floor_elevator1[21]), .out(n2003) );
  nand2 \eq_42_3/UGTI0_21  ( .a(n2002), .b(current_floor_output_elevator1[21]), 
        .out(\eq_42_3/GTV1 [21]) );
  nand2 \eq_42_3/UGTI1_21  ( .a(\eq_42_3/AEQB [21]), .b(\eq_42_3/GTV [21]), 
        .out(\eq_42_3/GTV2 [21]) );
  nand2 \eq_42_3/UGTI2_21  ( .a(\eq_42_3/GTV1 [21]), .b(\eq_42_3/GTV2 [21]), 
        .out(\eq_42_3/GTV [22]) );
  nand2 \eq_42_3/ULTI0_21  ( .a(n2001), .b(destination_floor_elevator1[21]), 
        .out(\eq_42_3/LTV1 [21]) );
  nand2 \eq_42_3/ULTI1_21  ( .a(\eq_42_3/AEQB [21]), .b(\eq_42_3/LTV [21]), 
        .out(\eq_42_3/LTV2 [21]) );
  nand2 \eq_42_3/ULTI2_21  ( .a(\eq_42_3/LTV1 [21]), .b(\eq_42_3/LTV2 [21]), 
        .out(\eq_42_3/LTV [22]) );
  xor2 \eq_42_3/UEQI_22  ( .a(current_floor_output_elevator1[22]), .b(
        destination_floor_elevator1[22]), .out(n2000) );
  nand2 \eq_42_3/UGTI0_22  ( .a(n1999), .b(current_floor_output_elevator1[22]), 
        .out(\eq_42_3/GTV1 [22]) );
  nand2 \eq_42_3/UGTI1_22  ( .a(\eq_42_3/AEQB [22]), .b(\eq_42_3/GTV [22]), 
        .out(\eq_42_3/GTV2 [22]) );
  nand2 \eq_42_3/UGTI2_22  ( .a(\eq_42_3/GTV1 [22]), .b(\eq_42_3/GTV2 [22]), 
        .out(\eq_42_3/GTV [23]) );
  nand2 \eq_42_3/ULTI0_22  ( .a(n1998), .b(destination_floor_elevator1[22]), 
        .out(\eq_42_3/LTV1 [22]) );
  nand2 \eq_42_3/ULTI1_22  ( .a(\eq_42_3/AEQB [22]), .b(\eq_42_3/LTV [22]), 
        .out(\eq_42_3/LTV2 [22]) );
  nand2 \eq_42_3/ULTI2_22  ( .a(\eq_42_3/LTV1 [22]), .b(\eq_42_3/LTV2 [22]), 
        .out(\eq_42_3/LTV [23]) );
  xor2 \eq_42_3/UEQI_23  ( .a(current_floor_output_elevator1[23]), .b(
        destination_floor_elevator1[23]), .out(n1997) );
  nand2 \eq_42_3/UGTI0_23  ( .a(n1996), .b(current_floor_output_elevator1[23]), 
        .out(\eq_42_3/GTV1 [23]) );
  nand2 \eq_42_3/UGTI1_23  ( .a(\eq_42_3/AEQB [23]), .b(\eq_42_3/GTV [23]), 
        .out(\eq_42_3/GTV2 [23]) );
  nand2 \eq_42_3/UGTI2_23  ( .a(\eq_42_3/GTV1 [23]), .b(\eq_42_3/GTV2 [23]), 
        .out(\eq_42_3/GTV [24]) );
  nand2 \eq_42_3/ULTI0_23  ( .a(n1995), .b(destination_floor_elevator1[23]), 
        .out(\eq_42_3/LTV1 [23]) );
  nand2 \eq_42_3/ULTI1_23  ( .a(\eq_42_3/AEQB [23]), .b(\eq_42_3/LTV [23]), 
        .out(\eq_42_3/LTV2 [23]) );
  nand2 \eq_42_3/ULTI2_23  ( .a(\eq_42_3/LTV1 [23]), .b(\eq_42_3/LTV2 [23]), 
        .out(\eq_42_3/LTV [24]) );
  xor2 \eq_42_3/UEQI_24  ( .a(current_floor_output_elevator1[24]), .b(
        destination_floor_elevator1[24]), .out(n1994) );
  nand2 \eq_42_3/UGTI0_24  ( .a(n1993), .b(current_floor_output_elevator1[24]), 
        .out(\eq_42_3/GTV1 [24]) );
  nand2 \eq_42_3/UGTI1_24  ( .a(\eq_42_3/AEQB [24]), .b(\eq_42_3/GTV [24]), 
        .out(\eq_42_3/GTV2 [24]) );
  nand2 \eq_42_3/UGTI2_24  ( .a(\eq_42_3/GTV1 [24]), .b(\eq_42_3/GTV2 [24]), 
        .out(\eq_42_3/GTV [25]) );
  nand2 \eq_42_3/ULTI0_24  ( .a(n1992), .b(destination_floor_elevator1[24]), 
        .out(\eq_42_3/LTV1 [24]) );
  nand2 \eq_42_3/ULTI1_24  ( .a(\eq_42_3/AEQB [24]), .b(\eq_42_3/LTV [24]), 
        .out(\eq_42_3/LTV2 [24]) );
  nand2 \eq_42_3/ULTI2_24  ( .a(\eq_42_3/LTV1 [24]), .b(\eq_42_3/LTV2 [24]), 
        .out(\eq_42_3/LTV [25]) );
  xor2 \eq_42_3/UEQI_25  ( .a(current_floor_output_elevator1[25]), .b(
        destination_floor_elevator1[25]), .out(n1991) );
  nand2 \eq_42_3/UGTI0_25  ( .a(n1990), .b(current_floor_output_elevator1[25]), 
        .out(\eq_42_3/GTV1 [25]) );
  nand2 \eq_42_3/UGTI1_25  ( .a(\eq_42_3/AEQB [25]), .b(\eq_42_3/GTV [25]), 
        .out(\eq_42_3/GTV2 [25]) );
  nand2 \eq_42_3/UGTI2_25  ( .a(\eq_42_3/GTV1 [25]), .b(\eq_42_3/GTV2 [25]), 
        .out(\eq_42_3/GTV [26]) );
  nand2 \eq_42_3/ULTI0_25  ( .a(n1989), .b(destination_floor_elevator1[25]), 
        .out(\eq_42_3/LTV1 [25]) );
  nand2 \eq_42_3/ULTI1_25  ( .a(\eq_42_3/AEQB [25]), .b(\eq_42_3/LTV [25]), 
        .out(\eq_42_3/LTV2 [25]) );
  nand2 \eq_42_3/ULTI2_25  ( .a(\eq_42_3/LTV1 [25]), .b(\eq_42_3/LTV2 [25]), 
        .out(\eq_42_3/LTV [26]) );
  xor2 \eq_42_3/UEQI_26  ( .a(current_floor_output_elevator1[26]), .b(
        destination_floor_elevator1[26]), .out(n1988) );
  nand2 \eq_42_3/UGTI0_26  ( .a(n1987), .b(current_floor_output_elevator1[26]), 
        .out(\eq_42_3/GTV1 [26]) );
  nand2 \eq_42_3/UGTI1_26  ( .a(\eq_42_3/AEQB [26]), .b(\eq_42_3/GTV [26]), 
        .out(\eq_42_3/GTV2 [26]) );
  nand2 \eq_42_3/UGTI2_26  ( .a(\eq_42_3/GTV1 [26]), .b(\eq_42_3/GTV2 [26]), 
        .out(\eq_42_3/GTV [27]) );
  nand2 \eq_42_3/ULTI0_26  ( .a(n1986), .b(destination_floor_elevator1[26]), 
        .out(\eq_42_3/LTV1 [26]) );
  nand2 \eq_42_3/ULTI1_26  ( .a(\eq_42_3/AEQB [26]), .b(\eq_42_3/LTV [26]), 
        .out(\eq_42_3/LTV2 [26]) );
  nand2 \eq_42_3/ULTI2_26  ( .a(\eq_42_3/LTV1 [26]), .b(\eq_42_3/LTV2 [26]), 
        .out(\eq_42_3/LTV [27]) );
  xor2 \eq_42_3/UEQI_27  ( .a(current_floor_output_elevator1[27]), .b(
        destination_floor_elevator1[27]), .out(n1985) );
  nand2 \eq_42_3/UGTI0_27  ( .a(n1984), .b(current_floor_output_elevator1[27]), 
        .out(\eq_42_3/GTV1 [27]) );
  nand2 \eq_42_3/UGTI1_27  ( .a(\eq_42_3/AEQB [27]), .b(\eq_42_3/GTV [27]), 
        .out(\eq_42_3/GTV2 [27]) );
  nand2 \eq_42_3/UGTI2_27  ( .a(\eq_42_3/GTV1 [27]), .b(\eq_42_3/GTV2 [27]), 
        .out(\eq_42_3/GTV [28]) );
  nand2 \eq_42_3/ULTI0_27  ( .a(n1983), .b(destination_floor_elevator1[27]), 
        .out(\eq_42_3/LTV1 [27]) );
  nand2 \eq_42_3/ULTI1_27  ( .a(\eq_42_3/AEQB [27]), .b(\eq_42_3/LTV [27]), 
        .out(\eq_42_3/LTV2 [27]) );
  nand2 \eq_42_3/ULTI2_27  ( .a(\eq_42_3/LTV1 [27]), .b(\eq_42_3/LTV2 [27]), 
        .out(\eq_42_3/LTV [28]) );
  xor2 \eq_42_3/UEQI_28  ( .a(current_floor_output_elevator1[28]), .b(
        destination_floor_elevator1[28]), .out(n1982) );
  nand2 \eq_42_3/UGTI0_28  ( .a(n1981), .b(current_floor_output_elevator1[28]), 
        .out(\eq_42_3/GTV1 [28]) );
  nand2 \eq_42_3/UGTI1_28  ( .a(\eq_42_3/AEQB [28]), .b(\eq_42_3/GTV [28]), 
        .out(\eq_42_3/GTV2 [28]) );
  nand2 \eq_42_3/UGTI2_28  ( .a(\eq_42_3/GTV1 [28]), .b(\eq_42_3/GTV2 [28]), 
        .out(\eq_42_3/GTV [29]) );
  nand2 \eq_42_3/ULTI0_28  ( .a(n1980), .b(destination_floor_elevator1[28]), 
        .out(\eq_42_3/LTV1 [28]) );
  nand2 \eq_42_3/ULTI1_28  ( .a(\eq_42_3/AEQB [28]), .b(\eq_42_3/LTV [28]), 
        .out(\eq_42_3/LTV2 [28]) );
  nand2 \eq_42_3/ULTI2_28  ( .a(\eq_42_3/LTV1 [28]), .b(\eq_42_3/LTV2 [28]), 
        .out(\eq_42_3/LTV [29]) );
  xor2 \eq_42_3/UEQI_29  ( .a(current_floor_output_elevator1[29]), .b(
        destination_floor_elevator1[29]), .out(n1979) );
  nand2 \eq_42_3/UGTI0_29  ( .a(n1978), .b(current_floor_output_elevator1[29]), 
        .out(\eq_42_3/GTV1 [29]) );
  nand2 \eq_42_3/UGTI1_29  ( .a(\eq_42_3/AEQB [29]), .b(\eq_42_3/GTV [29]), 
        .out(\eq_42_3/GTV2 [29]) );
  nand2 \eq_42_3/UGTI2_29  ( .a(\eq_42_3/GTV1 [29]), .b(\eq_42_3/GTV2 [29]), 
        .out(\eq_42_3/GTV [30]) );
  nand2 \eq_42_3/ULTI0_29  ( .a(n1977), .b(destination_floor_elevator1[29]), 
        .out(\eq_42_3/LTV1 [29]) );
  nand2 \eq_42_3/ULTI1_29  ( .a(\eq_42_3/AEQB [29]), .b(\eq_42_3/LTV [29]), 
        .out(\eq_42_3/LTV2 [29]) );
  nand2 \eq_42_3/ULTI2_29  ( .a(\eq_42_3/LTV1 [29]), .b(\eq_42_3/LTV2 [29]), 
        .out(\eq_42_3/LTV [30]) );
  xor2 \eq_42_3/UEQI_30  ( .a(current_floor_output_elevator1[30]), .b(
        destination_floor_elevator1[30]), .out(n1976) );
  nand2 \eq_42_3/UGTI0_30  ( .a(n1975), .b(current_floor_output_elevator1[30]), 
        .out(\eq_42_3/GTV1 [30]) );
  nand2 \eq_42_3/UGTI1_30  ( .a(\eq_42_3/AEQB [30]), .b(\eq_42_3/GTV [30]), 
        .out(\eq_42_3/GTV2 [30]) );
  nand2 \eq_42_3/UGTI2_30  ( .a(\eq_42_3/GTV1 [30]), .b(\eq_42_3/GTV2 [30]), 
        .out(\eq_42_3/GTV [31]) );
  nand2 \eq_42_3/ULTI0_30  ( .a(n1974), .b(destination_floor_elevator1[30]), 
        .out(\eq_42_3/LTV1 [30]) );
  nand2 \eq_42_3/ULTI1_30  ( .a(\eq_42_3/AEQB [30]), .b(\eq_42_3/LTV [30]), 
        .out(\eq_42_3/LTV2 [30]) );
  nand2 \eq_42_3/ULTI2_30  ( .a(\eq_42_3/LTV1 [30]), .b(\eq_42_3/LTV2 [30]), 
        .out(\eq_42_3/LTV [31]) );
  xor2 \eq_42_3/UEQI_31  ( .a(current_floor_output_elevator1[31]), .b(
        destination_floor_elevator1[31]), .out(n1973) );
  nand2 \eq_42_3/UGTI0_31  ( .a(n1972), .b(current_floor_output_elevator1[31]), 
        .out(\eq_42_3/GTV1 [31]) );
  nand2 \eq_42_3/UGTI1_31  ( .a(\eq_42_3/AEQB [31]), .b(\eq_42_3/GTV [31]), 
        .out(\eq_42_3/GTV2 [31]) );
  nand2 \eq_42_3/UGTI2_31  ( .a(\eq_42_3/GTV1 [31]), .b(\eq_42_3/GTV2 [31]), 
        .out(\eq_42_3/GTV [32]) );
  nand2 \eq_42_3/ULTI0_31  ( .a(n1971), .b(destination_floor_elevator1[31]), 
        .out(\eq_42_3/LTV1 [31]) );
  nand2 \eq_42_3/ULTI1_31  ( .a(\eq_42_3/AEQB [31]), .b(\eq_42_3/LTV [31]), 
        .out(\eq_42_3/LTV2 [31]) );
  nand2 \eq_42_3/ULTI2_31  ( .a(\eq_42_3/LTV1 [31]), .b(\eq_42_3/LTV2 [31]), 
        .out(\eq_42_3/LTV [32]) );
  xor2 \eq_42_3/UEQI_32  ( .a(current_floor_output_elevator1[32]), .b(
        destination_floor_elevator1[32]), .out(n1970) );
  nand2 \eq_42_3/UGTI0_32  ( .a(n1969), .b(current_floor_output_elevator1[32]), 
        .out(\eq_42_3/GTV1 [32]) );
  nand2 \eq_42_3/UGTI1_32  ( .a(\eq_42_3/AEQB [32]), .b(\eq_42_3/GTV [32]), 
        .out(\eq_42_3/GTV2 [32]) );
  nand2 \eq_42_3/UGTI2_32  ( .a(\eq_42_3/GTV1 [32]), .b(\eq_42_3/GTV2 [32]), 
        .out(\eq_42_3/GTV [33]) );
  nand2 \eq_42_3/ULTI0_32  ( .a(n1968), .b(destination_floor_elevator1[32]), 
        .out(\eq_42_3/LTV1 [32]) );
  nand2 \eq_42_3/ULTI1_32  ( .a(\eq_42_3/AEQB [32]), .b(\eq_42_3/LTV [32]), 
        .out(\eq_42_3/LTV2 [32]) );
  nand2 \eq_42_3/ULTI2_32  ( .a(\eq_42_3/LTV1 [32]), .b(\eq_42_3/LTV2 [32]), 
        .out(\eq_42_3/LTV [33]) );
  xor2 \eq_42_3/UEQI_33  ( .a(current_floor_output_elevator1[33]), .b(
        destination_floor_elevator1[33]), .out(n1967) );
  nand2 \eq_42_3/UGTI0_33  ( .a(n1966), .b(current_floor_output_elevator1[33]), 
        .out(\eq_42_3/GTV1 [33]) );
  nand2 \eq_42_3/UGTI1_33  ( .a(\eq_42_3/AEQB [33]), .b(\eq_42_3/GTV [33]), 
        .out(\eq_42_3/GTV2 [33]) );
  nand2 \eq_42_3/UGTI2_33  ( .a(\eq_42_3/GTV1 [33]), .b(\eq_42_3/GTV2 [33]), 
        .out(\eq_42_3/GTV [34]) );
  nand2 \eq_42_3/ULTI0_33  ( .a(n1965), .b(destination_floor_elevator1[33]), 
        .out(\eq_42_3/LTV1 [33]) );
  nand2 \eq_42_3/ULTI1_33  ( .a(\eq_42_3/AEQB [33]), .b(\eq_42_3/LTV [33]), 
        .out(\eq_42_3/LTV2 [33]) );
  nand2 \eq_42_3/ULTI2_33  ( .a(\eq_42_3/LTV1 [33]), .b(\eq_42_3/LTV2 [33]), 
        .out(\eq_42_3/LTV [34]) );
  xor2 \eq_42_3/UEQI_34  ( .a(current_floor_output_elevator1[34]), .b(
        destination_floor_elevator1[34]), .out(n1964) );
  nand2 \eq_42_3/UGTI0_34  ( .a(n1963), .b(current_floor_output_elevator1[34]), 
        .out(\eq_42_3/GTV1 [34]) );
  nand2 \eq_42_3/UGTI1_34  ( .a(\eq_42_3/AEQB [34]), .b(\eq_42_3/GTV [34]), 
        .out(\eq_42_3/GTV2 [34]) );
  nand2 \eq_42_3/UGTI2_34  ( .a(\eq_42_3/GTV1 [34]), .b(\eq_42_3/GTV2 [34]), 
        .out(\eq_42_3/GTV [35]) );
  nand2 \eq_42_3/ULTI0_34  ( .a(n1962), .b(destination_floor_elevator1[34]), 
        .out(\eq_42_3/LTV1 [34]) );
  nand2 \eq_42_3/ULTI1_34  ( .a(\eq_42_3/AEQB [34]), .b(\eq_42_3/LTV [34]), 
        .out(\eq_42_3/LTV2 [34]) );
  nand2 \eq_42_3/ULTI2_34  ( .a(\eq_42_3/LTV1 [34]), .b(\eq_42_3/LTV2 [34]), 
        .out(\eq_42_3/LTV [35]) );
  xor2 \eq_42_3/UEQI_35  ( .a(current_floor_output_elevator1[35]), .b(
        destination_floor_elevator1[35]), .out(n1961) );
  nand2 \eq_42_3/UGTI0_35  ( .a(n1960), .b(current_floor_output_elevator1[35]), 
        .out(\eq_42_3/GTV1 [35]) );
  nand2 \eq_42_3/UGTI1_35  ( .a(\eq_42_3/AEQB [35]), .b(\eq_42_3/GTV [35]), 
        .out(\eq_42_3/GTV2 [35]) );
  nand2 \eq_42_3/UGTI2_35  ( .a(\eq_42_3/GTV1 [35]), .b(\eq_42_3/GTV2 [35]), 
        .out(\eq_42_3/GTV [36]) );
  nand2 \eq_42_3/ULTI0_35  ( .a(n1959), .b(destination_floor_elevator1[35]), 
        .out(\eq_42_3/LTV1 [35]) );
  nand2 \eq_42_3/ULTI1_35  ( .a(\eq_42_3/AEQB [35]), .b(\eq_42_3/LTV [35]), 
        .out(\eq_42_3/LTV2 [35]) );
  nand2 \eq_42_3/ULTI2_35  ( .a(\eq_42_3/LTV1 [35]), .b(\eq_42_3/LTV2 [35]), 
        .out(\eq_42_3/LTV [36]) );
  xor2 \eq_42_3/UEQI_36  ( .a(current_floor_output_elevator1[36]), .b(
        destination_floor_elevator1[36]), .out(n1958) );
  nand2 \eq_42_3/UGTI0_36  ( .a(n1957), .b(current_floor_output_elevator1[36]), 
        .out(\eq_42_3/GTV1 [36]) );
  nand2 \eq_42_3/UGTI1_36  ( .a(\eq_42_3/AEQB [36]), .b(\eq_42_3/GTV [36]), 
        .out(\eq_42_3/GTV2 [36]) );
  nand2 \eq_42_3/UGTI2_36  ( .a(\eq_42_3/GTV1 [36]), .b(\eq_42_3/GTV2 [36]), 
        .out(\eq_42_3/GTV [37]) );
  nand2 \eq_42_3/ULTI0_36  ( .a(n1956), .b(destination_floor_elevator1[36]), 
        .out(\eq_42_3/LTV1 [36]) );
  nand2 \eq_42_3/ULTI1_36  ( .a(\eq_42_3/AEQB [36]), .b(\eq_42_3/LTV [36]), 
        .out(\eq_42_3/LTV2 [36]) );
  nand2 \eq_42_3/ULTI2_36  ( .a(\eq_42_3/LTV1 [36]), .b(\eq_42_3/LTV2 [36]), 
        .out(\eq_42_3/LTV [37]) );
  xor2 \eq_42_3/UEQI_37  ( .a(current_floor_output_elevator1[37]), .b(
        destination_floor_elevator1[37]), .out(n1955) );
  nand2 \eq_42_3/UGTI0_37  ( .a(n1954), .b(current_floor_output_elevator1[37]), 
        .out(\eq_42_3/GTV1 [37]) );
  nand2 \eq_42_3/UGTI1_37  ( .a(\eq_42_3/AEQB [37]), .b(\eq_42_3/GTV [37]), 
        .out(\eq_42_3/GTV2 [37]) );
  nand2 \eq_42_3/UGTI2_37  ( .a(\eq_42_3/GTV1 [37]), .b(\eq_42_3/GTV2 [37]), 
        .out(\eq_42_3/GTV [38]) );
  nand2 \eq_42_3/ULTI0_37  ( .a(n1953), .b(destination_floor_elevator1[37]), 
        .out(\eq_42_3/LTV1 [37]) );
  nand2 \eq_42_3/ULTI1_37  ( .a(\eq_42_3/AEQB [37]), .b(\eq_42_3/LTV [37]), 
        .out(\eq_42_3/LTV2 [37]) );
  nand2 \eq_42_3/ULTI2_37  ( .a(\eq_42_3/LTV1 [37]), .b(\eq_42_3/LTV2 [37]), 
        .out(\eq_42_3/LTV [38]) );
  xor2 \eq_42_3/UEQI_38  ( .a(current_floor_output_elevator1[38]), .b(
        destination_floor_elevator1[38]), .out(n1952) );
  nand2 \eq_42_3/UGTI0_38  ( .a(n1951), .b(current_floor_output_elevator1[38]), 
        .out(\eq_42_3/GTV1 [38]) );
  nand2 \eq_42_3/UGTI1_38  ( .a(\eq_42_3/AEQB [38]), .b(\eq_42_3/GTV [38]), 
        .out(\eq_42_3/GTV2 [38]) );
  nand2 \eq_42_3/UGTI2_38  ( .a(\eq_42_3/GTV1 [38]), .b(\eq_42_3/GTV2 [38]), 
        .out(\eq_42_3/GTV [39]) );
  nand2 \eq_42_3/ULTI0_38  ( .a(n1950), .b(destination_floor_elevator1[38]), 
        .out(\eq_42_3/LTV1 [38]) );
  nand2 \eq_42_3/ULTI1_38  ( .a(\eq_42_3/AEQB [38]), .b(\eq_42_3/LTV [38]), 
        .out(\eq_42_3/LTV2 [38]) );
  nand2 \eq_42_3/ULTI2_38  ( .a(\eq_42_3/LTV1 [38]), .b(\eq_42_3/LTV2 [38]), 
        .out(\eq_42_3/LTV [39]) );
  xor2 \eq_42_3/UEQI_39  ( .a(current_floor_output_elevator1[39]), .b(
        destination_floor_elevator1[39]), .out(n1949) );
  nand2 \eq_42_3/UGTI0_39  ( .a(n1948), .b(current_floor_output_elevator1[39]), 
        .out(\eq_42_3/GTV1 [39]) );
  nand2 \eq_42_3/UGTI1_39  ( .a(\eq_42_3/AEQB [39]), .b(\eq_42_3/GTV [39]), 
        .out(\eq_42_3/GTV2 [39]) );
  nand2 \eq_42_3/UGTI2_39  ( .a(\eq_42_3/GTV1 [39]), .b(\eq_42_3/GTV2 [39]), 
        .out(\eq_42_3/GTV [40]) );
  nand2 \eq_42_3/ULTI0_39  ( .a(n1947), .b(destination_floor_elevator1[39]), 
        .out(\eq_42_3/LTV1 [39]) );
  nand2 \eq_42_3/ULTI1_39  ( .a(\eq_42_3/AEQB [39]), .b(\eq_42_3/LTV [39]), 
        .out(\eq_42_3/LTV2 [39]) );
  nand2 \eq_42_3/ULTI2_39  ( .a(\eq_42_3/LTV1 [39]), .b(\eq_42_3/LTV2 [39]), 
        .out(\eq_42_3/LTV [40]) );
  xor2 \eq_42_3/UEQI_40  ( .a(current_floor_output_elevator1[40]), .b(
        destination_floor_elevator1[40]), .out(n1946) );
  nand2 \eq_42_3/UGTI0_40  ( .a(n1945), .b(current_floor_output_elevator1[40]), 
        .out(\eq_42_3/GTV1 [40]) );
  nand2 \eq_42_3/UGTI1_40  ( .a(\eq_42_3/AEQB [40]), .b(\eq_42_3/GTV [40]), 
        .out(\eq_42_3/GTV2 [40]) );
  nand2 \eq_42_3/UGTI2_40  ( .a(\eq_42_3/GTV1 [40]), .b(\eq_42_3/GTV2 [40]), 
        .out(\eq_42_3/GTV [41]) );
  nand2 \eq_42_3/ULTI0_40  ( .a(n1944), .b(destination_floor_elevator1[40]), 
        .out(\eq_42_3/LTV1 [40]) );
  nand2 \eq_42_3/ULTI1_40  ( .a(\eq_42_3/AEQB [40]), .b(\eq_42_3/LTV [40]), 
        .out(\eq_42_3/LTV2 [40]) );
  nand2 \eq_42_3/ULTI2_40  ( .a(\eq_42_3/LTV1 [40]), .b(\eq_42_3/LTV2 [40]), 
        .out(\eq_42_3/LTV [41]) );
  xor2 \eq_42_3/UEQI_41  ( .a(current_floor_output_elevator1[41]), .b(
        destination_floor_elevator1[41]), .out(n1943) );
  nand2 \eq_42_3/UGTI0_41  ( .a(n1942), .b(current_floor_output_elevator1[41]), 
        .out(\eq_42_3/GTV1 [41]) );
  nand2 \eq_42_3/UGTI1_41  ( .a(\eq_42_3/AEQB [41]), .b(\eq_42_3/GTV [41]), 
        .out(\eq_42_3/GTV2 [41]) );
  nand2 \eq_42_3/UGTI2_41  ( .a(\eq_42_3/GTV1 [41]), .b(\eq_42_3/GTV2 [41]), 
        .out(\eq_42_3/GTV [42]) );
  nand2 \eq_42_3/ULTI0_41  ( .a(n1941), .b(destination_floor_elevator1[41]), 
        .out(\eq_42_3/LTV1 [41]) );
  nand2 \eq_42_3/ULTI1_41  ( .a(\eq_42_3/AEQB [41]), .b(\eq_42_3/LTV [41]), 
        .out(\eq_42_3/LTV2 [41]) );
  nand2 \eq_42_3/ULTI2_41  ( .a(\eq_42_3/LTV1 [41]), .b(\eq_42_3/LTV2 [41]), 
        .out(\eq_42_3/LTV [42]) );
  xor2 \eq_42_3/UEQI_42  ( .a(current_floor_output_elevator1[42]), .b(
        destination_floor_elevator1[42]), .out(n1940) );
  nand2 \eq_42_3/UGTI0_42  ( .a(n1939), .b(current_floor_output_elevator1[42]), 
        .out(\eq_42_3/GTV1 [42]) );
  nand2 \eq_42_3/UGTI1_42  ( .a(\eq_42_3/AEQB [42]), .b(\eq_42_3/GTV [42]), 
        .out(\eq_42_3/GTV2 [42]) );
  nand2 \eq_42_3/UGTI2_42  ( .a(\eq_42_3/GTV1 [42]), .b(\eq_42_3/GTV2 [42]), 
        .out(\eq_42_3/GTV [43]) );
  nand2 \eq_42_3/ULTI0_42  ( .a(n1938), .b(destination_floor_elevator1[42]), 
        .out(\eq_42_3/LTV1 [42]) );
  nand2 \eq_42_3/ULTI1_42  ( .a(\eq_42_3/AEQB [42]), .b(\eq_42_3/LTV [42]), 
        .out(\eq_42_3/LTV2 [42]) );
  nand2 \eq_42_3/ULTI2_42  ( .a(\eq_42_3/LTV1 [42]), .b(\eq_42_3/LTV2 [42]), 
        .out(\eq_42_3/LTV [43]) );
  xor2 \eq_42_3/UEQI_43  ( .a(current_floor_output_elevator1[43]), .b(
        destination_floor_elevator1[43]), .out(n1937) );
  nand2 \eq_42_3/UGTI0_43  ( .a(n1936), .b(current_floor_output_elevator1[43]), 
        .out(\eq_42_3/GTV1 [43]) );
  nand2 \eq_42_3/UGTI1_43  ( .a(\eq_42_3/AEQB [43]), .b(\eq_42_3/GTV [43]), 
        .out(\eq_42_3/GTV2 [43]) );
  nand2 \eq_42_3/UGTI2_43  ( .a(\eq_42_3/GTV1 [43]), .b(\eq_42_3/GTV2 [43]), 
        .out(\eq_42_3/GTV [44]) );
  nand2 \eq_42_3/ULTI0_43  ( .a(n1935), .b(destination_floor_elevator1[43]), 
        .out(\eq_42_3/LTV1 [43]) );
  nand2 \eq_42_3/ULTI1_43  ( .a(\eq_42_3/AEQB [43]), .b(\eq_42_3/LTV [43]), 
        .out(\eq_42_3/LTV2 [43]) );
  nand2 \eq_42_3/ULTI2_43  ( .a(\eq_42_3/LTV1 [43]), .b(\eq_42_3/LTV2 [43]), 
        .out(\eq_42_3/LTV [44]) );
  xor2 \eq_42_3/UEQI_44  ( .a(current_floor_output_elevator1[44]), .b(
        destination_floor_elevator1[44]), .out(n1934) );
  nand2 \eq_42_3/UGTI0_44  ( .a(n1933), .b(current_floor_output_elevator1[44]), 
        .out(\eq_42_3/GTV1 [44]) );
  nand2 \eq_42_3/UGTI1_44  ( .a(\eq_42_3/AEQB [44]), .b(\eq_42_3/GTV [44]), 
        .out(\eq_42_3/GTV2 [44]) );
  nand2 \eq_42_3/UGTI2_44  ( .a(\eq_42_3/GTV1 [44]), .b(\eq_42_3/GTV2 [44]), 
        .out(\eq_42_3/GTV [45]) );
  nand2 \eq_42_3/ULTI0_44  ( .a(n1932), .b(destination_floor_elevator1[44]), 
        .out(\eq_42_3/LTV1 [44]) );
  nand2 \eq_42_3/ULTI1_44  ( .a(\eq_42_3/AEQB [44]), .b(\eq_42_3/LTV [44]), 
        .out(\eq_42_3/LTV2 [44]) );
  nand2 \eq_42_3/ULTI2_44  ( .a(\eq_42_3/LTV1 [44]), .b(\eq_42_3/LTV2 [44]), 
        .out(\eq_42_3/LTV [45]) );
  xor2 \eq_42_3/UEQI_45  ( .a(current_floor_output_elevator1[45]), .b(
        destination_floor_elevator1[45]), .out(n1931) );
  nand2 \eq_42_3/UGTI0_45  ( .a(n1930), .b(current_floor_output_elevator1[45]), 
        .out(\eq_42_3/GTV1 [45]) );
  nand2 \eq_42_3/UGTI1_45  ( .a(\eq_42_3/AEQB [45]), .b(\eq_42_3/GTV [45]), 
        .out(\eq_42_3/GTV2 [45]) );
  nand2 \eq_42_3/UGTI2_45  ( .a(\eq_42_3/GTV1 [45]), .b(\eq_42_3/GTV2 [45]), 
        .out(\eq_42_3/GTV [46]) );
  nand2 \eq_42_3/ULTI0_45  ( .a(n1929), .b(destination_floor_elevator1[45]), 
        .out(\eq_42_3/LTV1 [45]) );
  nand2 \eq_42_3/ULTI1_45  ( .a(\eq_42_3/AEQB [45]), .b(\eq_42_3/LTV [45]), 
        .out(\eq_42_3/LTV2 [45]) );
  nand2 \eq_42_3/ULTI2_45  ( .a(\eq_42_3/LTV1 [45]), .b(\eq_42_3/LTV2 [45]), 
        .out(\eq_42_3/LTV [46]) );
  xor2 \eq_42_3/UEQI_46  ( .a(current_floor_output_elevator1[46]), .b(
        destination_floor_elevator1[46]), .out(n1928) );
  nand2 \eq_42_3/UGTI0_46  ( .a(n1927), .b(current_floor_output_elevator1[46]), 
        .out(\eq_42_3/GTV1 [46]) );
  nand2 \eq_42_3/UGTI1_46  ( .a(\eq_42_3/AEQB [46]), .b(\eq_42_3/GTV [46]), 
        .out(\eq_42_3/GTV2 [46]) );
  nand2 \eq_42_3/UGTI2_46  ( .a(\eq_42_3/GTV1 [46]), .b(\eq_42_3/GTV2 [46]), 
        .out(\eq_42_3/GTV [47]) );
  nand2 \eq_42_3/ULTI0_46  ( .a(n1926), .b(destination_floor_elevator1[46]), 
        .out(\eq_42_3/LTV1 [46]) );
  nand2 \eq_42_3/ULTI1_46  ( .a(\eq_42_3/AEQB [46]), .b(\eq_42_3/LTV [46]), 
        .out(\eq_42_3/LTV2 [46]) );
  nand2 \eq_42_3/ULTI2_46  ( .a(\eq_42_3/LTV1 [46]), .b(\eq_42_3/LTV2 [46]), 
        .out(\eq_42_3/LTV [47]) );
  xor2 \eq_42_3/UEQI_47  ( .a(current_floor_output_elevator1[47]), .b(
        destination_floor_elevator1[47]), .out(n1925) );
  nand2 \eq_42_3/UGTI0_47  ( .a(n1924), .b(current_floor_output_elevator1[47]), 
        .out(\eq_42_3/GTV1 [47]) );
  nand2 \eq_42_3/UGTI1_47  ( .a(\eq_42_3/AEQB [47]), .b(\eq_42_3/GTV [47]), 
        .out(\eq_42_3/GTV2 [47]) );
  nand2 \eq_42_3/UGTI2_47  ( .a(\eq_42_3/GTV1 [47]), .b(\eq_42_3/GTV2 [47]), 
        .out(\eq_42_3/GTV [48]) );
  nand2 \eq_42_3/ULTI0_47  ( .a(n1923), .b(destination_floor_elevator1[47]), 
        .out(\eq_42_3/LTV1 [47]) );
  nand2 \eq_42_3/ULTI1_47  ( .a(\eq_42_3/AEQB [47]), .b(\eq_42_3/LTV [47]), 
        .out(\eq_42_3/LTV2 [47]) );
  nand2 \eq_42_3/ULTI2_47  ( .a(\eq_42_3/LTV1 [47]), .b(\eq_42_3/LTV2 [47]), 
        .out(\eq_42_3/LTV [48]) );
  xor2 \eq_42_3/UEQI_48  ( .a(current_floor_output_elevator1[48]), .b(
        destination_floor_elevator1[48]), .out(n1922) );
  nand2 \eq_42_3/UGTI0_48  ( .a(n1921), .b(current_floor_output_elevator1[48]), 
        .out(\eq_42_3/GTV1 [48]) );
  nand2 \eq_42_3/UGTI1_48  ( .a(\eq_42_3/AEQB [48]), .b(\eq_42_3/GTV [48]), 
        .out(\eq_42_3/GTV2 [48]) );
  nand2 \eq_42_3/UGTI2_48  ( .a(\eq_42_3/GTV1 [48]), .b(\eq_42_3/GTV2 [48]), 
        .out(\eq_42_3/GTV [49]) );
  nand2 \eq_42_3/ULTI0_48  ( .a(n1920), .b(destination_floor_elevator1[48]), 
        .out(\eq_42_3/LTV1 [48]) );
  nand2 \eq_42_3/ULTI1_48  ( .a(\eq_42_3/AEQB [48]), .b(\eq_42_3/LTV [48]), 
        .out(\eq_42_3/LTV2 [48]) );
  nand2 \eq_42_3/ULTI2_48  ( .a(\eq_42_3/LTV1 [48]), .b(\eq_42_3/LTV2 [48]), 
        .out(\eq_42_3/LTV [49]) );
  xor2 \eq_42_3/UEQI_49  ( .a(current_floor_output_elevator1[49]), .b(
        destination_floor_elevator1[49]), .out(n1919) );
  nand2 \eq_42_3/UGTI0_49  ( .a(n1918), .b(current_floor_output_elevator1[49]), 
        .out(\eq_42_3/GTV1 [49]) );
  nand2 \eq_42_3/UGTI1_49  ( .a(\eq_42_3/AEQB [49]), .b(\eq_42_3/GTV [49]), 
        .out(\eq_42_3/GTV2 [49]) );
  nand2 \eq_42_3/UGTI2_49  ( .a(\eq_42_3/GTV1 [49]), .b(\eq_42_3/GTV2 [49]), 
        .out(\eq_42_3/GTV [50]) );
  nand2 \eq_42_3/ULTI0_49  ( .a(n1917), .b(destination_floor_elevator1[49]), 
        .out(\eq_42_3/LTV1 [49]) );
  nand2 \eq_42_3/ULTI1_49  ( .a(\eq_42_3/AEQB [49]), .b(\eq_42_3/LTV [49]), 
        .out(\eq_42_3/LTV2 [49]) );
  nand2 \eq_42_3/ULTI2_49  ( .a(\eq_42_3/LTV1 [49]), .b(\eq_42_3/LTV2 [49]), 
        .out(\eq_42_3/LTV [50]) );
  xor2 \eq_42_3/UEQI_50  ( .a(current_floor_output_elevator1[50]), .b(
        destination_floor_elevator1[50]), .out(n1916) );
  nand2 \eq_42_3/UGTI0_50  ( .a(n1915), .b(current_floor_output_elevator1[50]), 
        .out(\eq_42_3/GTV1 [50]) );
  nand2 \eq_42_3/UGTI1_50  ( .a(\eq_42_3/AEQB [50]), .b(\eq_42_3/GTV [50]), 
        .out(\eq_42_3/GTV2 [50]) );
  nand2 \eq_42_3/UGTI2_50  ( .a(\eq_42_3/GTV1 [50]), .b(\eq_42_3/GTV2 [50]), 
        .out(\eq_42_3/GTV [51]) );
  nand2 \eq_42_3/ULTI0_50  ( .a(n1914), .b(destination_floor_elevator1[50]), 
        .out(\eq_42_3/LTV1 [50]) );
  nand2 \eq_42_3/ULTI1_50  ( .a(\eq_42_3/AEQB [50]), .b(\eq_42_3/LTV [50]), 
        .out(\eq_42_3/LTV2 [50]) );
  nand2 \eq_42_3/ULTI2_50  ( .a(\eq_42_3/LTV1 [50]), .b(\eq_42_3/LTV2 [50]), 
        .out(\eq_42_3/LTV [51]) );
  xor2 \eq_42_3/UEQI_51  ( .a(current_floor_output_elevator1[51]), .b(
        destination_floor_elevator1[51]), .out(n1913) );
  nand2 \eq_42_3/UGTI0_51  ( .a(n1912), .b(current_floor_output_elevator1[51]), 
        .out(\eq_42_3/GTV1 [51]) );
  nand2 \eq_42_3/UGTI1_51  ( .a(\eq_42_3/AEQB [51]), .b(\eq_42_3/GTV [51]), 
        .out(\eq_42_3/GTV2 [51]) );
  nand2 \eq_42_3/UGTI2_51  ( .a(\eq_42_3/GTV1 [51]), .b(\eq_42_3/GTV2 [51]), 
        .out(\eq_42_3/GTV [52]) );
  nand2 \eq_42_3/ULTI0_51  ( .a(n1911), .b(destination_floor_elevator1[51]), 
        .out(\eq_42_3/LTV1 [51]) );
  nand2 \eq_42_3/ULTI1_51  ( .a(\eq_42_3/AEQB [51]), .b(\eq_42_3/LTV [51]), 
        .out(\eq_42_3/LTV2 [51]) );
  nand2 \eq_42_3/ULTI2_51  ( .a(\eq_42_3/LTV1 [51]), .b(\eq_42_3/LTV2 [51]), 
        .out(\eq_42_3/LTV [52]) );
  xor2 \eq_42_3/UEQI_52  ( .a(current_floor_output_elevator1[52]), .b(
        destination_floor_elevator1[52]), .out(n1910) );
  nand2 \eq_42_3/UGTI0_52  ( .a(n1909), .b(current_floor_output_elevator1[52]), 
        .out(\eq_42_3/GTV1 [52]) );
  nand2 \eq_42_3/UGTI1_52  ( .a(\eq_42_3/AEQB [52]), .b(\eq_42_3/GTV [52]), 
        .out(\eq_42_3/GTV2 [52]) );
  nand2 \eq_42_3/UGTI2_52  ( .a(\eq_42_3/GTV1 [52]), .b(\eq_42_3/GTV2 [52]), 
        .out(\eq_42_3/GTV [53]) );
  nand2 \eq_42_3/ULTI0_52  ( .a(n1908), .b(destination_floor_elevator1[52]), 
        .out(\eq_42_3/LTV1 [52]) );
  nand2 \eq_42_3/ULTI1_52  ( .a(\eq_42_3/AEQB [52]), .b(\eq_42_3/LTV [52]), 
        .out(\eq_42_3/LTV2 [52]) );
  nand2 \eq_42_3/ULTI2_52  ( .a(\eq_42_3/LTV1 [52]), .b(\eq_42_3/LTV2 [52]), 
        .out(\eq_42_3/LTV [53]) );
  xor2 \eq_42_3/UEQI_53  ( .a(current_floor_output_elevator1[53]), .b(
        destination_floor_elevator1[53]), .out(n1907) );
  nand2 \eq_42_3/UGTI0_53  ( .a(n1906), .b(current_floor_output_elevator1[53]), 
        .out(\eq_42_3/GTV1 [53]) );
  nand2 \eq_42_3/UGTI1_53  ( .a(\eq_42_3/AEQB [53]), .b(\eq_42_3/GTV [53]), 
        .out(\eq_42_3/GTV2 [53]) );
  nand2 \eq_42_3/UGTI2_53  ( .a(\eq_42_3/GTV1 [53]), .b(\eq_42_3/GTV2 [53]), 
        .out(\eq_42_3/GTV [54]) );
  nand2 \eq_42_3/ULTI0_53  ( .a(n1905), .b(destination_floor_elevator1[53]), 
        .out(\eq_42_3/LTV1 [53]) );
  nand2 \eq_42_3/ULTI1_53  ( .a(\eq_42_3/AEQB [53]), .b(\eq_42_3/LTV [53]), 
        .out(\eq_42_3/LTV2 [53]) );
  nand2 \eq_42_3/ULTI2_53  ( .a(\eq_42_3/LTV1 [53]), .b(\eq_42_3/LTV2 [53]), 
        .out(\eq_42_3/LTV [54]) );
  xor2 \eq_42_3/UEQI_54  ( .a(current_floor_output_elevator1[54]), .b(
        destination_floor_elevator1[54]), .out(n1904) );
  nand2 \eq_42_3/UGTI0_54  ( .a(n1903), .b(current_floor_output_elevator1[54]), 
        .out(\eq_42_3/GTV1 [54]) );
  nand2 \eq_42_3/UGTI1_54  ( .a(\eq_42_3/AEQB [54]), .b(\eq_42_3/GTV [54]), 
        .out(\eq_42_3/GTV2 [54]) );
  nand2 \eq_42_3/UGTI2_54  ( .a(\eq_42_3/GTV1 [54]), .b(\eq_42_3/GTV2 [54]), 
        .out(\eq_42_3/GTV [55]) );
  nand2 \eq_42_3/ULTI0_54  ( .a(n1902), .b(destination_floor_elevator1[54]), 
        .out(\eq_42_3/LTV1 [54]) );
  nand2 \eq_42_3/ULTI1_54  ( .a(\eq_42_3/AEQB [54]), .b(\eq_42_3/LTV [54]), 
        .out(\eq_42_3/LTV2 [54]) );
  nand2 \eq_42_3/ULTI2_54  ( .a(\eq_42_3/LTV1 [54]), .b(\eq_42_3/LTV2 [54]), 
        .out(\eq_42_3/LTV [55]) );
  xor2 \eq_42_3/UEQI_55  ( .a(current_floor_output_elevator1[55]), .b(
        destination_floor_elevator1[55]), .out(n1901) );
  nand2 \eq_42_3/UGTI0_55  ( .a(n1900), .b(current_floor_output_elevator1[55]), 
        .out(\eq_42_3/GTV1 [55]) );
  nand2 \eq_42_3/UGTI1_55  ( .a(\eq_42_3/AEQB [55]), .b(\eq_42_3/GTV [55]), 
        .out(\eq_42_3/GTV2 [55]) );
  nand2 \eq_42_3/UGTI2_55  ( .a(\eq_42_3/GTV1 [55]), .b(\eq_42_3/GTV2 [55]), 
        .out(\eq_42_3/GTV [56]) );
  nand2 \eq_42_3/ULTI0_55  ( .a(n1899), .b(destination_floor_elevator1[55]), 
        .out(\eq_42_3/LTV1 [55]) );
  nand2 \eq_42_3/ULTI1_55  ( .a(\eq_42_3/AEQB [55]), .b(\eq_42_3/LTV [55]), 
        .out(\eq_42_3/LTV2 [55]) );
  nand2 \eq_42_3/ULTI2_55  ( .a(\eq_42_3/LTV1 [55]), .b(\eq_42_3/LTV2 [55]), 
        .out(\eq_42_3/LTV [56]) );
  xor2 \eq_42_3/UEQI_56  ( .a(current_floor_output_elevator1[56]), .b(
        destination_floor_elevator1[56]), .out(n1898) );
  nand2 \eq_42_3/UGTI0_56  ( .a(n1897), .b(current_floor_output_elevator1[56]), 
        .out(\eq_42_3/GTV1 [56]) );
  nand2 \eq_42_3/UGTI1_56  ( .a(\eq_42_3/AEQB [56]), .b(\eq_42_3/GTV [56]), 
        .out(\eq_42_3/GTV2 [56]) );
  nand2 \eq_42_3/UGTI2_56  ( .a(\eq_42_3/GTV1 [56]), .b(\eq_42_3/GTV2 [56]), 
        .out(\eq_42_3/GTV [57]) );
  nand2 \eq_42_3/ULTI0_56  ( .a(n1896), .b(destination_floor_elevator1[56]), 
        .out(\eq_42_3/LTV1 [56]) );
  nand2 \eq_42_3/ULTI1_56  ( .a(\eq_42_3/AEQB [56]), .b(\eq_42_3/LTV [56]), 
        .out(\eq_42_3/LTV2 [56]) );
  nand2 \eq_42_3/ULTI2_56  ( .a(\eq_42_3/LTV1 [56]), .b(\eq_42_3/LTV2 [56]), 
        .out(\eq_42_3/LTV [57]) );
  xor2 \eq_42_3/UEQI_57  ( .a(current_floor_output_elevator1[57]), .b(
        destination_floor_elevator1[57]), .out(n1895) );
  nand2 \eq_42_3/UGTI0_57  ( .a(n1894), .b(current_floor_output_elevator1[57]), 
        .out(\eq_42_3/GTV1 [57]) );
  nand2 \eq_42_3/UGTI1_57  ( .a(\eq_42_3/AEQB [57]), .b(\eq_42_3/GTV [57]), 
        .out(\eq_42_3/GTV2 [57]) );
  nand2 \eq_42_3/UGTI2_57  ( .a(\eq_42_3/GTV1 [57]), .b(\eq_42_3/GTV2 [57]), 
        .out(\eq_42_3/GTV [58]) );
  nand2 \eq_42_3/ULTI0_57  ( .a(n1893), .b(destination_floor_elevator1[57]), 
        .out(\eq_42_3/LTV1 [57]) );
  nand2 \eq_42_3/ULTI1_57  ( .a(\eq_42_3/AEQB [57]), .b(\eq_42_3/LTV [57]), 
        .out(\eq_42_3/LTV2 [57]) );
  nand2 \eq_42_3/ULTI2_57  ( .a(\eq_42_3/LTV1 [57]), .b(\eq_42_3/LTV2 [57]), 
        .out(\eq_42_3/LTV [58]) );
  xor2 \eq_42_3/UEQI_58  ( .a(current_floor_output_elevator1[58]), .b(
        destination_floor_elevator1[58]), .out(n1892) );
  nand2 \eq_42_3/UGTI0_58  ( .a(n1891), .b(current_floor_output_elevator1[58]), 
        .out(\eq_42_3/GTV1 [58]) );
  nand2 \eq_42_3/UGTI1_58  ( .a(\eq_42_3/AEQB [58]), .b(\eq_42_3/GTV [58]), 
        .out(\eq_42_3/GTV2 [58]) );
  nand2 \eq_42_3/UGTI2_58  ( .a(\eq_42_3/GTV1 [58]), .b(\eq_42_3/GTV2 [58]), 
        .out(\eq_42_3/GTV [59]) );
  nand2 \eq_42_3/ULTI0_58  ( .a(n1890), .b(destination_floor_elevator1[58]), 
        .out(\eq_42_3/LTV1 [58]) );
  nand2 \eq_42_3/ULTI1_58  ( .a(\eq_42_3/AEQB [58]), .b(\eq_42_3/LTV [58]), 
        .out(\eq_42_3/LTV2 [58]) );
  nand2 \eq_42_3/ULTI2_58  ( .a(\eq_42_3/LTV1 [58]), .b(\eq_42_3/LTV2 [58]), 
        .out(\eq_42_3/LTV [59]) );
  xor2 \eq_42_3/UEQI_59  ( .a(current_floor_output_elevator1[59]), .b(
        destination_floor_elevator1[59]), .out(n1889) );
  nand2 \eq_42_3/UGTI0_59  ( .a(n1888), .b(current_floor_output_elevator1[59]), 
        .out(\eq_42_3/GTV1 [59]) );
  nand2 \eq_42_3/UGTI1_59  ( .a(\eq_42_3/AEQB [59]), .b(\eq_42_3/GTV [59]), 
        .out(\eq_42_3/GTV2 [59]) );
  nand2 \eq_42_3/UGTI2_59  ( .a(\eq_42_3/GTV1 [59]), .b(\eq_42_3/GTV2 [59]), 
        .out(\eq_42_3/GTV [60]) );
  nand2 \eq_42_3/ULTI0_59  ( .a(n1887), .b(destination_floor_elevator1[59]), 
        .out(\eq_42_3/LTV1 [59]) );
  nand2 \eq_42_3/ULTI1_59  ( .a(\eq_42_3/AEQB [59]), .b(\eq_42_3/LTV [59]), 
        .out(\eq_42_3/LTV2 [59]) );
  nand2 \eq_42_3/ULTI2_59  ( .a(\eq_42_3/LTV1 [59]), .b(\eq_42_3/LTV2 [59]), 
        .out(\eq_42_3/LTV [60]) );
  xor2 \eq_42_3/UEQI_60  ( .a(current_floor_output_elevator1[60]), .b(
        destination_floor_elevator1[60]), .out(n1886) );
  nand2 \eq_42_3/UGTI0_60  ( .a(n1885), .b(current_floor_output_elevator1[60]), 
        .out(\eq_42_3/GTV1 [60]) );
  nand2 \eq_42_3/UGTI1_60  ( .a(\eq_42_3/AEQB [60]), .b(\eq_42_3/GTV [60]), 
        .out(\eq_42_3/GTV2 [60]) );
  nand2 \eq_42_3/UGTI2_60  ( .a(\eq_42_3/GTV1 [60]), .b(\eq_42_3/GTV2 [60]), 
        .out(\eq_42_3/GTV [61]) );
  nand2 \eq_42_3/ULTI0_60  ( .a(n1884), .b(destination_floor_elevator1[60]), 
        .out(\eq_42_3/LTV1 [60]) );
  nand2 \eq_42_3/ULTI1_60  ( .a(\eq_42_3/AEQB [60]), .b(\eq_42_3/LTV [60]), 
        .out(\eq_42_3/LTV2 [60]) );
  nand2 \eq_42_3/ULTI2_60  ( .a(\eq_42_3/LTV1 [60]), .b(\eq_42_3/LTV2 [60]), 
        .out(\eq_42_3/LTV [61]) );
  xor2 \eq_42_3/UEQI_61  ( .a(current_floor_output_elevator1[61]), .b(
        destination_floor_elevator1[61]), .out(n1883) );
  nand2 \eq_42_3/UGTI0_61  ( .a(n1882), .b(current_floor_output_elevator1[61]), 
        .out(\eq_42_3/GTV1 [61]) );
  nand2 \eq_42_3/UGTI1_61  ( .a(\eq_42_3/AEQB [61]), .b(\eq_42_3/GTV [61]), 
        .out(\eq_42_3/GTV2 [61]) );
  nand2 \eq_42_3/UGTI2_61  ( .a(\eq_42_3/GTV1 [61]), .b(\eq_42_3/GTV2 [61]), 
        .out(\eq_42_3/GTV [62]) );
  nand2 \eq_42_3/ULTI0_61  ( .a(n1881), .b(destination_floor_elevator1[61]), 
        .out(\eq_42_3/LTV1 [61]) );
  nand2 \eq_42_3/ULTI1_61  ( .a(\eq_42_3/AEQB [61]), .b(\eq_42_3/LTV [61]), 
        .out(\eq_42_3/LTV2 [61]) );
  nand2 \eq_42_3/ULTI2_61  ( .a(\eq_42_3/LTV1 [61]), .b(\eq_42_3/LTV2 [61]), 
        .out(\eq_42_3/LTV [62]) );
  xor2 \eq_42_3/UEQI_62  ( .a(current_floor_output_elevator1[62]), .b(
        destination_floor_elevator1[62]), .out(n1880) );
  nand2 \eq_42_3/UGTI0_62  ( .a(n1879), .b(current_floor_output_elevator1[62]), 
        .out(\eq_42_3/GTV1 [62]) );
  nand2 \eq_42_3/UGTI1_62  ( .a(\eq_42_3/AEQB [62]), .b(\eq_42_3/GTV [62]), 
        .out(\eq_42_3/GTV2 [62]) );
  nand2 \eq_42_3/UGTI2_62  ( .a(\eq_42_3/GTV1 [62]), .b(\eq_42_3/GTV2 [62]), 
        .out(\eq_42_3/GTV [63]) );
  nand2 \eq_42_3/ULTI0_62  ( .a(n1878), .b(destination_floor_elevator1[62]), 
        .out(\eq_42_3/LTV1 [62]) );
  nand2 \eq_42_3/ULTI1_62  ( .a(\eq_42_3/AEQB [62]), .b(\eq_42_3/LTV [62]), 
        .out(\eq_42_3/LTV2 [62]) );
  nand2 \eq_42_3/ULTI2_62  ( .a(\eq_42_3/LTV1 [62]), .b(\eq_42_3/LTV2 [62]), 
        .out(\eq_42_3/LTV [63]) );
  nor2 \ne_42/UEQ  ( .a(\ne_42/GT ), .b(\ne_42/LT ), .out(\ne_42/EQ ) );
  inv \ne_42/UNE  ( .in(\ne_42/EQ ), .out(N12) );
  nand2 \ne_42/UNGT0  ( .a(final_floor_elevator2[0]), .b(n1877), .out(n1876)
         );
  nand2 \ne_42/UNLT0  ( .a(requested_floor[0]), .b(n1875), .out(n1874) );
  xor2 \ne_42/UEQI  ( .a(\ne_42/SA ), .b(\ne_47/SB ), .out(n1873) );
  nand2 \ne_42/UGTI0  ( .a(n1872), .b(\ne_42/SA ), .out(\ne_42/GTV1 [63]) );
  nand2 \ne_42/UGTI1  ( .a(\ne_42/AEQB [63]), .b(\ne_42/GTV [63]), .out(
        \ne_42/GTV2 [63]) );
  nand2 \ne_42/UGTI2  ( .a(\ne_42/GTV1 [63]), .b(\ne_42/GTV2 [63]), .out(
        \ne_42/GT ) );
  nand2 \ne_42/ULTI0  ( .a(n1871), .b(\ne_47/SB ), .out(\ne_42/LTV1 [63]) );
  nand2 \ne_42/ULTI1  ( .a(\ne_42/AEQB [63]), .b(\ne_42/LTV [63]), .out(
        \ne_42/LTV2 [63]) );
  nand2 \ne_42/ULTI2  ( .a(\ne_42/LTV1 [63]), .b(\ne_42/LTV2 [63]), .out(
        \ne_42/LT ) );
  xor2 \ne_42/UEQI_1  ( .a(final_floor_elevator2[1]), .b(requested_floor[1]), 
        .out(n1870) );
  nand2 \ne_42/UGTI0_1  ( .a(n1869), .b(final_floor_elevator2[1]), .out(
        \ne_42/GTV1 [1]) );
  nand2 \ne_42/UGTI1_1  ( .a(\ne_42/AEQB [1]), .b(\ne_42/GTV [1]), .out(
        \ne_42/GTV2 [1]) );
  nand2 \ne_42/UGTI2_1  ( .a(\ne_42/GTV1 [1]), .b(\ne_42/GTV2 [1]), .out(
        \ne_42/GTV [2]) );
  nand2 \ne_42/ULTI0_1  ( .a(n1868), .b(requested_floor[1]), .out(
        \ne_42/LTV1 [1]) );
  nand2 \ne_42/ULTI1_1  ( .a(\ne_42/AEQB [1]), .b(\ne_42/LTV [1]), .out(
        \ne_42/LTV2 [1]) );
  nand2 \ne_42/ULTI2_1  ( .a(\ne_42/LTV1 [1]), .b(\ne_42/LTV2 [1]), .out(
        \ne_42/LTV [2]) );
  xor2 \ne_42/UEQI_2  ( .a(final_floor_elevator2[2]), .b(requested_floor[2]), 
        .out(n1867) );
  nand2 \ne_42/UGTI0_2  ( .a(n1866), .b(final_floor_elevator2[2]), .out(
        \ne_42/GTV1 [2]) );
  nand2 \ne_42/UGTI1_2  ( .a(\ne_42/AEQB [2]), .b(\ne_42/GTV [2]), .out(
        \ne_42/GTV2 [2]) );
  nand2 \ne_42/UGTI2_2  ( .a(\ne_42/GTV1 [2]), .b(\ne_42/GTV2 [2]), .out(
        \ne_42/GTV [3]) );
  nand2 \ne_42/ULTI0_2  ( .a(n1865), .b(requested_floor[2]), .out(
        \ne_42/LTV1 [2]) );
  nand2 \ne_42/ULTI1_2  ( .a(\ne_42/AEQB [2]), .b(\ne_42/LTV [2]), .out(
        \ne_42/LTV2 [2]) );
  nand2 \ne_42/ULTI2_2  ( .a(\ne_42/LTV1 [2]), .b(\ne_42/LTV2 [2]), .out(
        \ne_42/LTV [3]) );
  xor2 \ne_42/UEQI_3  ( .a(final_floor_elevator2[3]), .b(requested_floor[3]), 
        .out(n1864) );
  nand2 \ne_42/UGTI0_3  ( .a(n1863), .b(final_floor_elevator2[3]), .out(
        \ne_42/GTV1 [3]) );
  nand2 \ne_42/UGTI1_3  ( .a(\ne_42/AEQB [3]), .b(\ne_42/GTV [3]), .out(
        \ne_42/GTV2 [3]) );
  nand2 \ne_42/UGTI2_3  ( .a(\ne_42/GTV1 [3]), .b(\ne_42/GTV2 [3]), .out(
        \ne_42/GTV [4]) );
  nand2 \ne_42/ULTI0_3  ( .a(n1862), .b(requested_floor[3]), .out(
        \ne_42/LTV1 [3]) );
  nand2 \ne_42/ULTI1_3  ( .a(\ne_42/AEQB [3]), .b(\ne_42/LTV [3]), .out(
        \ne_42/LTV2 [3]) );
  nand2 \ne_42/ULTI2_3  ( .a(\ne_42/LTV1 [3]), .b(\ne_42/LTV2 [3]), .out(
        \ne_42/LTV [4]) );
  xor2 \ne_42/UEQI_4  ( .a(final_floor_elevator2[4]), .b(requested_floor[4]), 
        .out(n1861) );
  nand2 \ne_42/UGTI0_4  ( .a(n1860), .b(final_floor_elevator2[4]), .out(
        \ne_42/GTV1 [4]) );
  nand2 \ne_42/UGTI1_4  ( .a(\ne_42/AEQB [4]), .b(\ne_42/GTV [4]), .out(
        \ne_42/GTV2 [4]) );
  nand2 \ne_42/UGTI2_4  ( .a(\ne_42/GTV1 [4]), .b(\ne_42/GTV2 [4]), .out(
        \ne_42/GTV [5]) );
  nand2 \ne_42/ULTI0_4  ( .a(n1859), .b(requested_floor[4]), .out(
        \ne_42/LTV1 [4]) );
  nand2 \ne_42/ULTI1_4  ( .a(\ne_42/AEQB [4]), .b(\ne_42/LTV [4]), .out(
        \ne_42/LTV2 [4]) );
  nand2 \ne_42/ULTI2_4  ( .a(\ne_42/LTV1 [4]), .b(\ne_42/LTV2 [4]), .out(
        \ne_42/LTV [5]) );
  xor2 \ne_42/UEQI_5  ( .a(final_floor_elevator2[5]), .b(requested_floor[5]), 
        .out(n1858) );
  nand2 \ne_42/UGTI0_5  ( .a(n1857), .b(final_floor_elevator2[5]), .out(
        \ne_42/GTV1 [5]) );
  nand2 \ne_42/UGTI1_5  ( .a(\ne_42/AEQB [5]), .b(\ne_42/GTV [5]), .out(
        \ne_42/GTV2 [5]) );
  nand2 \ne_42/UGTI2_5  ( .a(\ne_42/GTV1 [5]), .b(\ne_42/GTV2 [5]), .out(
        \ne_42/GTV [6]) );
  nand2 \ne_42/ULTI0_5  ( .a(n1856), .b(requested_floor[5]), .out(
        \ne_42/LTV1 [5]) );
  nand2 \ne_42/ULTI1_5  ( .a(\ne_42/AEQB [5]), .b(\ne_42/LTV [5]), .out(
        \ne_42/LTV2 [5]) );
  nand2 \ne_42/ULTI2_5  ( .a(\ne_42/LTV1 [5]), .b(\ne_42/LTV2 [5]), .out(
        \ne_42/LTV [6]) );
  xor2 \ne_42/UEQI_6  ( .a(final_floor_elevator2[6]), .b(requested_floor[6]), 
        .out(n1855) );
  nand2 \ne_42/UGTI0_6  ( .a(n1854), .b(final_floor_elevator2[6]), .out(
        \ne_42/GTV1 [6]) );
  nand2 \ne_42/UGTI1_6  ( .a(\ne_42/AEQB [6]), .b(\ne_42/GTV [6]), .out(
        \ne_42/GTV2 [6]) );
  nand2 \ne_42/UGTI2_6  ( .a(\ne_42/GTV1 [6]), .b(\ne_42/GTV2 [6]), .out(
        \ne_42/GTV [7]) );
  nand2 \ne_42/ULTI0_6  ( .a(n1853), .b(requested_floor[6]), .out(
        \ne_42/LTV1 [6]) );
  nand2 \ne_42/ULTI1_6  ( .a(\ne_42/AEQB [6]), .b(\ne_42/LTV [6]), .out(
        \ne_42/LTV2 [6]) );
  nand2 \ne_42/ULTI2_6  ( .a(\ne_42/LTV1 [6]), .b(\ne_42/LTV2 [6]), .out(
        \ne_42/LTV [7]) );
  xor2 \ne_42/UEQI_7  ( .a(final_floor_elevator2[7]), .b(requested_floor[7]), 
        .out(n1852) );
  nand2 \ne_42/UGTI0_7  ( .a(n1851), .b(final_floor_elevator2[7]), .out(
        \ne_42/GTV1 [7]) );
  nand2 \ne_42/UGTI1_7  ( .a(\ne_42/AEQB [7]), .b(\ne_42/GTV [7]), .out(
        \ne_42/GTV2 [7]) );
  nand2 \ne_42/UGTI2_7  ( .a(\ne_42/GTV1 [7]), .b(\ne_42/GTV2 [7]), .out(
        \ne_42/GTV [8]) );
  nand2 \ne_42/ULTI0_7  ( .a(n1850), .b(requested_floor[7]), .out(
        \ne_42/LTV1 [7]) );
  nand2 \ne_42/ULTI1_7  ( .a(\ne_42/AEQB [7]), .b(\ne_42/LTV [7]), .out(
        \ne_42/LTV2 [7]) );
  nand2 \ne_42/ULTI2_7  ( .a(\ne_42/LTV1 [7]), .b(\ne_42/LTV2 [7]), .out(
        \ne_42/LTV [8]) );
  xor2 \ne_42/UEQI_8  ( .a(final_floor_elevator2[8]), .b(requested_floor[8]), 
        .out(n1849) );
  nand2 \ne_42/UGTI0_8  ( .a(n1848), .b(final_floor_elevator2[8]), .out(
        \ne_42/GTV1 [8]) );
  nand2 \ne_42/UGTI1_8  ( .a(\ne_42/AEQB [8]), .b(\ne_42/GTV [8]), .out(
        \ne_42/GTV2 [8]) );
  nand2 \ne_42/UGTI2_8  ( .a(\ne_42/GTV1 [8]), .b(\ne_42/GTV2 [8]), .out(
        \ne_42/GTV [9]) );
  nand2 \ne_42/ULTI0_8  ( .a(n1847), .b(requested_floor[8]), .out(
        \ne_42/LTV1 [8]) );
  nand2 \ne_42/ULTI1_8  ( .a(\ne_42/AEQB [8]), .b(\ne_42/LTV [8]), .out(
        \ne_42/LTV2 [8]) );
  nand2 \ne_42/ULTI2_8  ( .a(\ne_42/LTV1 [8]), .b(\ne_42/LTV2 [8]), .out(
        \ne_42/LTV [9]) );
  xor2 \ne_42/UEQI_9  ( .a(final_floor_elevator2[9]), .b(requested_floor[9]), 
        .out(n1846) );
  nand2 \ne_42/UGTI0_9  ( .a(n1845), .b(final_floor_elevator2[9]), .out(
        \ne_42/GTV1 [9]) );
  nand2 \ne_42/UGTI1_9  ( .a(\ne_42/AEQB [9]), .b(\ne_42/GTV [9]), .out(
        \ne_42/GTV2 [9]) );
  nand2 \ne_42/UGTI2_9  ( .a(\ne_42/GTV1 [9]), .b(\ne_42/GTV2 [9]), .out(
        \ne_42/GTV [10]) );
  nand2 \ne_42/ULTI0_9  ( .a(n1844), .b(requested_floor[9]), .out(
        \ne_42/LTV1 [9]) );
  nand2 \ne_42/ULTI1_9  ( .a(\ne_42/AEQB [9]), .b(\ne_42/LTV [9]), .out(
        \ne_42/LTV2 [9]) );
  nand2 \ne_42/ULTI2_9  ( .a(\ne_42/LTV1 [9]), .b(\ne_42/LTV2 [9]), .out(
        \ne_42/LTV [10]) );
  xor2 \ne_42/UEQI_10  ( .a(final_floor_elevator2[10]), .b(requested_floor[10]), .out(n1843) );
  nand2 \ne_42/UGTI0_10  ( .a(n1842), .b(final_floor_elevator2[10]), .out(
        \ne_42/GTV1 [10]) );
  nand2 \ne_42/UGTI1_10  ( .a(\ne_42/AEQB [10]), .b(\ne_42/GTV [10]), .out(
        \ne_42/GTV2 [10]) );
  nand2 \ne_42/UGTI2_10  ( .a(\ne_42/GTV1 [10]), .b(\ne_42/GTV2 [10]), .out(
        \ne_42/GTV [11]) );
  nand2 \ne_42/ULTI0_10  ( .a(n1841), .b(requested_floor[10]), .out(
        \ne_42/LTV1 [10]) );
  nand2 \ne_42/ULTI1_10  ( .a(\ne_42/AEQB [10]), .b(\ne_42/LTV [10]), .out(
        \ne_42/LTV2 [10]) );
  nand2 \ne_42/ULTI2_10  ( .a(\ne_42/LTV1 [10]), .b(\ne_42/LTV2 [10]), .out(
        \ne_42/LTV [11]) );
  xor2 \ne_42/UEQI_11  ( .a(final_floor_elevator2[11]), .b(requested_floor[11]), .out(n1840) );
  nand2 \ne_42/UGTI0_11  ( .a(n1839), .b(final_floor_elevator2[11]), .out(
        \ne_42/GTV1 [11]) );
  nand2 \ne_42/UGTI1_11  ( .a(\ne_42/AEQB [11]), .b(\ne_42/GTV [11]), .out(
        \ne_42/GTV2 [11]) );
  nand2 \ne_42/UGTI2_11  ( .a(\ne_42/GTV1 [11]), .b(\ne_42/GTV2 [11]), .out(
        \ne_42/GTV [12]) );
  nand2 \ne_42/ULTI0_11  ( .a(n1838), .b(requested_floor[11]), .out(
        \ne_42/LTV1 [11]) );
  nand2 \ne_42/ULTI1_11  ( .a(\ne_42/AEQB [11]), .b(\ne_42/LTV [11]), .out(
        \ne_42/LTV2 [11]) );
  nand2 \ne_42/ULTI2_11  ( .a(\ne_42/LTV1 [11]), .b(\ne_42/LTV2 [11]), .out(
        \ne_42/LTV [12]) );
  xor2 \ne_42/UEQI_12  ( .a(final_floor_elevator2[12]), .b(requested_floor[12]), .out(n1837) );
  nand2 \ne_42/UGTI0_12  ( .a(n1836), .b(final_floor_elevator2[12]), .out(
        \ne_42/GTV1 [12]) );
  nand2 \ne_42/UGTI1_12  ( .a(\ne_42/AEQB [12]), .b(\ne_42/GTV [12]), .out(
        \ne_42/GTV2 [12]) );
  nand2 \ne_42/UGTI2_12  ( .a(\ne_42/GTV1 [12]), .b(\ne_42/GTV2 [12]), .out(
        \ne_42/GTV [13]) );
  nand2 \ne_42/ULTI0_12  ( .a(n1835), .b(requested_floor[12]), .out(
        \ne_42/LTV1 [12]) );
  nand2 \ne_42/ULTI1_12  ( .a(\ne_42/AEQB [12]), .b(\ne_42/LTV [12]), .out(
        \ne_42/LTV2 [12]) );
  nand2 \ne_42/ULTI2_12  ( .a(\ne_42/LTV1 [12]), .b(\ne_42/LTV2 [12]), .out(
        \ne_42/LTV [13]) );
  xor2 \ne_42/UEQI_13  ( .a(final_floor_elevator2[13]), .b(requested_floor[13]), .out(n1834) );
  nand2 \ne_42/UGTI0_13  ( .a(n1833), .b(final_floor_elevator2[13]), .out(
        \ne_42/GTV1 [13]) );
  nand2 \ne_42/UGTI1_13  ( .a(\ne_42/AEQB [13]), .b(\ne_42/GTV [13]), .out(
        \ne_42/GTV2 [13]) );
  nand2 \ne_42/UGTI2_13  ( .a(\ne_42/GTV1 [13]), .b(\ne_42/GTV2 [13]), .out(
        \ne_42/GTV [14]) );
  nand2 \ne_42/ULTI0_13  ( .a(n1832), .b(requested_floor[13]), .out(
        \ne_42/LTV1 [13]) );
  nand2 \ne_42/ULTI1_13  ( .a(\ne_42/AEQB [13]), .b(\ne_42/LTV [13]), .out(
        \ne_42/LTV2 [13]) );
  nand2 \ne_42/ULTI2_13  ( .a(\ne_42/LTV1 [13]), .b(\ne_42/LTV2 [13]), .out(
        \ne_42/LTV [14]) );
  xor2 \ne_42/UEQI_14  ( .a(final_floor_elevator2[14]), .b(requested_floor[14]), .out(n1831) );
  nand2 \ne_42/UGTI0_14  ( .a(n1830), .b(final_floor_elevator2[14]), .out(
        \ne_42/GTV1 [14]) );
  nand2 \ne_42/UGTI1_14  ( .a(\ne_42/AEQB [14]), .b(\ne_42/GTV [14]), .out(
        \ne_42/GTV2 [14]) );
  nand2 \ne_42/UGTI2_14  ( .a(\ne_42/GTV1 [14]), .b(\ne_42/GTV2 [14]), .out(
        \ne_42/GTV [15]) );
  nand2 \ne_42/ULTI0_14  ( .a(n1829), .b(requested_floor[14]), .out(
        \ne_42/LTV1 [14]) );
  nand2 \ne_42/ULTI1_14  ( .a(\ne_42/AEQB [14]), .b(\ne_42/LTV [14]), .out(
        \ne_42/LTV2 [14]) );
  nand2 \ne_42/ULTI2_14  ( .a(\ne_42/LTV1 [14]), .b(\ne_42/LTV2 [14]), .out(
        \ne_42/LTV [15]) );
  xor2 \ne_42/UEQI_15  ( .a(final_floor_elevator2[15]), .b(requested_floor[15]), .out(n1828) );
  nand2 \ne_42/UGTI0_15  ( .a(n1827), .b(final_floor_elevator2[15]), .out(
        \ne_42/GTV1 [15]) );
  nand2 \ne_42/UGTI1_15  ( .a(\ne_42/AEQB [15]), .b(\ne_42/GTV [15]), .out(
        \ne_42/GTV2 [15]) );
  nand2 \ne_42/UGTI2_15  ( .a(\ne_42/GTV1 [15]), .b(\ne_42/GTV2 [15]), .out(
        \ne_42/GTV [16]) );
  nand2 \ne_42/ULTI0_15  ( .a(n1826), .b(requested_floor[15]), .out(
        \ne_42/LTV1 [15]) );
  nand2 \ne_42/ULTI1_15  ( .a(\ne_42/AEQB [15]), .b(\ne_42/LTV [15]), .out(
        \ne_42/LTV2 [15]) );
  nand2 \ne_42/ULTI2_15  ( .a(\ne_42/LTV1 [15]), .b(\ne_42/LTV2 [15]), .out(
        \ne_42/LTV [16]) );
  xor2 \ne_42/UEQI_16  ( .a(final_floor_elevator2[16]), .b(requested_floor[16]), .out(n1825) );
  nand2 \ne_42/UGTI0_16  ( .a(n1824), .b(final_floor_elevator2[16]), .out(
        \ne_42/GTV1 [16]) );
  nand2 \ne_42/UGTI1_16  ( .a(\ne_42/AEQB [16]), .b(\ne_42/GTV [16]), .out(
        \ne_42/GTV2 [16]) );
  nand2 \ne_42/UGTI2_16  ( .a(\ne_42/GTV1 [16]), .b(\ne_42/GTV2 [16]), .out(
        \ne_42/GTV [17]) );
  nand2 \ne_42/ULTI0_16  ( .a(n1823), .b(requested_floor[16]), .out(
        \ne_42/LTV1 [16]) );
  nand2 \ne_42/ULTI1_16  ( .a(\ne_42/AEQB [16]), .b(\ne_42/LTV [16]), .out(
        \ne_42/LTV2 [16]) );
  nand2 \ne_42/ULTI2_16  ( .a(\ne_42/LTV1 [16]), .b(\ne_42/LTV2 [16]), .out(
        \ne_42/LTV [17]) );
  xor2 \ne_42/UEQI_17  ( .a(final_floor_elevator2[17]), .b(requested_floor[17]), .out(n1822) );
  nand2 \ne_42/UGTI0_17  ( .a(n1821), .b(final_floor_elevator2[17]), .out(
        \ne_42/GTV1 [17]) );
  nand2 \ne_42/UGTI1_17  ( .a(\ne_42/AEQB [17]), .b(\ne_42/GTV [17]), .out(
        \ne_42/GTV2 [17]) );
  nand2 \ne_42/UGTI2_17  ( .a(\ne_42/GTV1 [17]), .b(\ne_42/GTV2 [17]), .out(
        \ne_42/GTV [18]) );
  nand2 \ne_42/ULTI0_17  ( .a(n1820), .b(requested_floor[17]), .out(
        \ne_42/LTV1 [17]) );
  nand2 \ne_42/ULTI1_17  ( .a(\ne_42/AEQB [17]), .b(\ne_42/LTV [17]), .out(
        \ne_42/LTV2 [17]) );
  nand2 \ne_42/ULTI2_17  ( .a(\ne_42/LTV1 [17]), .b(\ne_42/LTV2 [17]), .out(
        \ne_42/LTV [18]) );
  xor2 \ne_42/UEQI_18  ( .a(final_floor_elevator2[18]), .b(requested_floor[18]), .out(n1819) );
  nand2 \ne_42/UGTI0_18  ( .a(n1818), .b(final_floor_elevator2[18]), .out(
        \ne_42/GTV1 [18]) );
  nand2 \ne_42/UGTI1_18  ( .a(\ne_42/AEQB [18]), .b(\ne_42/GTV [18]), .out(
        \ne_42/GTV2 [18]) );
  nand2 \ne_42/UGTI2_18  ( .a(\ne_42/GTV1 [18]), .b(\ne_42/GTV2 [18]), .out(
        \ne_42/GTV [19]) );
  nand2 \ne_42/ULTI0_18  ( .a(n1817), .b(requested_floor[18]), .out(
        \ne_42/LTV1 [18]) );
  nand2 \ne_42/ULTI1_18  ( .a(\ne_42/AEQB [18]), .b(\ne_42/LTV [18]), .out(
        \ne_42/LTV2 [18]) );
  nand2 \ne_42/ULTI2_18  ( .a(\ne_42/LTV1 [18]), .b(\ne_42/LTV2 [18]), .out(
        \ne_42/LTV [19]) );
  xor2 \ne_42/UEQI_19  ( .a(final_floor_elevator2[19]), .b(requested_floor[19]), .out(n1816) );
  nand2 \ne_42/UGTI0_19  ( .a(n1815), .b(final_floor_elevator2[19]), .out(
        \ne_42/GTV1 [19]) );
  nand2 \ne_42/UGTI1_19  ( .a(\ne_42/AEQB [19]), .b(\ne_42/GTV [19]), .out(
        \ne_42/GTV2 [19]) );
  nand2 \ne_42/UGTI2_19  ( .a(\ne_42/GTV1 [19]), .b(\ne_42/GTV2 [19]), .out(
        \ne_42/GTV [20]) );
  nand2 \ne_42/ULTI0_19  ( .a(n1814), .b(requested_floor[19]), .out(
        \ne_42/LTV1 [19]) );
  nand2 \ne_42/ULTI1_19  ( .a(\ne_42/AEQB [19]), .b(\ne_42/LTV [19]), .out(
        \ne_42/LTV2 [19]) );
  nand2 \ne_42/ULTI2_19  ( .a(\ne_42/LTV1 [19]), .b(\ne_42/LTV2 [19]), .out(
        \ne_42/LTV [20]) );
  xor2 \ne_42/UEQI_20  ( .a(final_floor_elevator2[20]), .b(requested_floor[20]), .out(n1813) );
  nand2 \ne_42/UGTI0_20  ( .a(n1812), .b(final_floor_elevator2[20]), .out(
        \ne_42/GTV1 [20]) );
  nand2 \ne_42/UGTI1_20  ( .a(\ne_42/AEQB [20]), .b(\ne_42/GTV [20]), .out(
        \ne_42/GTV2 [20]) );
  nand2 \ne_42/UGTI2_20  ( .a(\ne_42/GTV1 [20]), .b(\ne_42/GTV2 [20]), .out(
        \ne_42/GTV [21]) );
  nand2 \ne_42/ULTI0_20  ( .a(n1811), .b(requested_floor[20]), .out(
        \ne_42/LTV1 [20]) );
  nand2 \ne_42/ULTI1_20  ( .a(\ne_42/AEQB [20]), .b(\ne_42/LTV [20]), .out(
        \ne_42/LTV2 [20]) );
  nand2 \ne_42/ULTI2_20  ( .a(\ne_42/LTV1 [20]), .b(\ne_42/LTV2 [20]), .out(
        \ne_42/LTV [21]) );
  xor2 \ne_42/UEQI_21  ( .a(final_floor_elevator2[21]), .b(requested_floor[21]), .out(n1810) );
  nand2 \ne_42/UGTI0_21  ( .a(n1809), .b(final_floor_elevator2[21]), .out(
        \ne_42/GTV1 [21]) );
  nand2 \ne_42/UGTI1_21  ( .a(\ne_42/AEQB [21]), .b(\ne_42/GTV [21]), .out(
        \ne_42/GTV2 [21]) );
  nand2 \ne_42/UGTI2_21  ( .a(\ne_42/GTV1 [21]), .b(\ne_42/GTV2 [21]), .out(
        \ne_42/GTV [22]) );
  nand2 \ne_42/ULTI0_21  ( .a(n1808), .b(requested_floor[21]), .out(
        \ne_42/LTV1 [21]) );
  nand2 \ne_42/ULTI1_21  ( .a(\ne_42/AEQB [21]), .b(\ne_42/LTV [21]), .out(
        \ne_42/LTV2 [21]) );
  nand2 \ne_42/ULTI2_21  ( .a(\ne_42/LTV1 [21]), .b(\ne_42/LTV2 [21]), .out(
        \ne_42/LTV [22]) );
  xor2 \ne_42/UEQI_22  ( .a(final_floor_elevator2[22]), .b(requested_floor[22]), .out(n1807) );
  nand2 \ne_42/UGTI0_22  ( .a(n1806), .b(final_floor_elevator2[22]), .out(
        \ne_42/GTV1 [22]) );
  nand2 \ne_42/UGTI1_22  ( .a(\ne_42/AEQB [22]), .b(\ne_42/GTV [22]), .out(
        \ne_42/GTV2 [22]) );
  nand2 \ne_42/UGTI2_22  ( .a(\ne_42/GTV1 [22]), .b(\ne_42/GTV2 [22]), .out(
        \ne_42/GTV [23]) );
  nand2 \ne_42/ULTI0_22  ( .a(n1805), .b(requested_floor[22]), .out(
        \ne_42/LTV1 [22]) );
  nand2 \ne_42/ULTI1_22  ( .a(\ne_42/AEQB [22]), .b(\ne_42/LTV [22]), .out(
        \ne_42/LTV2 [22]) );
  nand2 \ne_42/ULTI2_22  ( .a(\ne_42/LTV1 [22]), .b(\ne_42/LTV2 [22]), .out(
        \ne_42/LTV [23]) );
  xor2 \ne_42/UEQI_23  ( .a(final_floor_elevator2[23]), .b(requested_floor[23]), .out(n1804) );
  nand2 \ne_42/UGTI0_23  ( .a(n1803), .b(final_floor_elevator2[23]), .out(
        \ne_42/GTV1 [23]) );
  nand2 \ne_42/UGTI1_23  ( .a(\ne_42/AEQB [23]), .b(\ne_42/GTV [23]), .out(
        \ne_42/GTV2 [23]) );
  nand2 \ne_42/UGTI2_23  ( .a(\ne_42/GTV1 [23]), .b(\ne_42/GTV2 [23]), .out(
        \ne_42/GTV [24]) );
  nand2 \ne_42/ULTI0_23  ( .a(n1802), .b(requested_floor[23]), .out(
        \ne_42/LTV1 [23]) );
  nand2 \ne_42/ULTI1_23  ( .a(\ne_42/AEQB [23]), .b(\ne_42/LTV [23]), .out(
        \ne_42/LTV2 [23]) );
  nand2 \ne_42/ULTI2_23  ( .a(\ne_42/LTV1 [23]), .b(\ne_42/LTV2 [23]), .out(
        \ne_42/LTV [24]) );
  xor2 \ne_42/UEQI_24  ( .a(final_floor_elevator2[24]), .b(requested_floor[24]), .out(n1801) );
  nand2 \ne_42/UGTI0_24  ( .a(n1800), .b(final_floor_elevator2[24]), .out(
        \ne_42/GTV1 [24]) );
  nand2 \ne_42/UGTI1_24  ( .a(\ne_42/AEQB [24]), .b(\ne_42/GTV [24]), .out(
        \ne_42/GTV2 [24]) );
  nand2 \ne_42/UGTI2_24  ( .a(\ne_42/GTV1 [24]), .b(\ne_42/GTV2 [24]), .out(
        \ne_42/GTV [25]) );
  nand2 \ne_42/ULTI0_24  ( .a(n1799), .b(requested_floor[24]), .out(
        \ne_42/LTV1 [24]) );
  nand2 \ne_42/ULTI1_24  ( .a(\ne_42/AEQB [24]), .b(\ne_42/LTV [24]), .out(
        \ne_42/LTV2 [24]) );
  nand2 \ne_42/ULTI2_24  ( .a(\ne_42/LTV1 [24]), .b(\ne_42/LTV2 [24]), .out(
        \ne_42/LTV [25]) );
  xor2 \ne_42/UEQI_25  ( .a(final_floor_elevator2[25]), .b(requested_floor[25]), .out(n1798) );
  nand2 \ne_42/UGTI0_25  ( .a(n1797), .b(final_floor_elevator2[25]), .out(
        \ne_42/GTV1 [25]) );
  nand2 \ne_42/UGTI1_25  ( .a(\ne_42/AEQB [25]), .b(\ne_42/GTV [25]), .out(
        \ne_42/GTV2 [25]) );
  nand2 \ne_42/UGTI2_25  ( .a(\ne_42/GTV1 [25]), .b(\ne_42/GTV2 [25]), .out(
        \ne_42/GTV [26]) );
  nand2 \ne_42/ULTI0_25  ( .a(n1796), .b(requested_floor[25]), .out(
        \ne_42/LTV1 [25]) );
  nand2 \ne_42/ULTI1_25  ( .a(\ne_42/AEQB [25]), .b(\ne_42/LTV [25]), .out(
        \ne_42/LTV2 [25]) );
  nand2 \ne_42/ULTI2_25  ( .a(\ne_42/LTV1 [25]), .b(\ne_42/LTV2 [25]), .out(
        \ne_42/LTV [26]) );
  xor2 \ne_42/UEQI_26  ( .a(final_floor_elevator2[26]), .b(requested_floor[26]), .out(n1795) );
  nand2 \ne_42/UGTI0_26  ( .a(n1794), .b(final_floor_elevator2[26]), .out(
        \ne_42/GTV1 [26]) );
  nand2 \ne_42/UGTI1_26  ( .a(\ne_42/AEQB [26]), .b(\ne_42/GTV [26]), .out(
        \ne_42/GTV2 [26]) );
  nand2 \ne_42/UGTI2_26  ( .a(\ne_42/GTV1 [26]), .b(\ne_42/GTV2 [26]), .out(
        \ne_42/GTV [27]) );
  nand2 \ne_42/ULTI0_26  ( .a(n1793), .b(requested_floor[26]), .out(
        \ne_42/LTV1 [26]) );
  nand2 \ne_42/ULTI1_26  ( .a(\ne_42/AEQB [26]), .b(\ne_42/LTV [26]), .out(
        \ne_42/LTV2 [26]) );
  nand2 \ne_42/ULTI2_26  ( .a(\ne_42/LTV1 [26]), .b(\ne_42/LTV2 [26]), .out(
        \ne_42/LTV [27]) );
  xor2 \ne_42/UEQI_27  ( .a(final_floor_elevator2[27]), .b(requested_floor[27]), .out(n1792) );
  nand2 \ne_42/UGTI0_27  ( .a(n1791), .b(final_floor_elevator2[27]), .out(
        \ne_42/GTV1 [27]) );
  nand2 \ne_42/UGTI1_27  ( .a(\ne_42/AEQB [27]), .b(\ne_42/GTV [27]), .out(
        \ne_42/GTV2 [27]) );
  nand2 \ne_42/UGTI2_27  ( .a(\ne_42/GTV1 [27]), .b(\ne_42/GTV2 [27]), .out(
        \ne_42/GTV [28]) );
  nand2 \ne_42/ULTI0_27  ( .a(n1790), .b(requested_floor[27]), .out(
        \ne_42/LTV1 [27]) );
  nand2 \ne_42/ULTI1_27  ( .a(\ne_42/AEQB [27]), .b(\ne_42/LTV [27]), .out(
        \ne_42/LTV2 [27]) );
  nand2 \ne_42/ULTI2_27  ( .a(\ne_42/LTV1 [27]), .b(\ne_42/LTV2 [27]), .out(
        \ne_42/LTV [28]) );
  xor2 \ne_42/UEQI_28  ( .a(final_floor_elevator2[28]), .b(requested_floor[28]), .out(n1789) );
  nand2 \ne_42/UGTI0_28  ( .a(n1788), .b(final_floor_elevator2[28]), .out(
        \ne_42/GTV1 [28]) );
  nand2 \ne_42/UGTI1_28  ( .a(\ne_42/AEQB [28]), .b(\ne_42/GTV [28]), .out(
        \ne_42/GTV2 [28]) );
  nand2 \ne_42/UGTI2_28  ( .a(\ne_42/GTV1 [28]), .b(\ne_42/GTV2 [28]), .out(
        \ne_42/GTV [29]) );
  nand2 \ne_42/ULTI0_28  ( .a(n1787), .b(requested_floor[28]), .out(
        \ne_42/LTV1 [28]) );
  nand2 \ne_42/ULTI1_28  ( .a(\ne_42/AEQB [28]), .b(\ne_42/LTV [28]), .out(
        \ne_42/LTV2 [28]) );
  nand2 \ne_42/ULTI2_28  ( .a(\ne_42/LTV1 [28]), .b(\ne_42/LTV2 [28]), .out(
        \ne_42/LTV [29]) );
  xor2 \ne_42/UEQI_29  ( .a(final_floor_elevator2[29]), .b(requested_floor[29]), .out(n1786) );
  nand2 \ne_42/UGTI0_29  ( .a(n1785), .b(final_floor_elevator2[29]), .out(
        \ne_42/GTV1 [29]) );
  nand2 \ne_42/UGTI1_29  ( .a(\ne_42/AEQB [29]), .b(\ne_42/GTV [29]), .out(
        \ne_42/GTV2 [29]) );
  nand2 \ne_42/UGTI2_29  ( .a(\ne_42/GTV1 [29]), .b(\ne_42/GTV2 [29]), .out(
        \ne_42/GTV [30]) );
  nand2 \ne_42/ULTI0_29  ( .a(n1784), .b(requested_floor[29]), .out(
        \ne_42/LTV1 [29]) );
  nand2 \ne_42/ULTI1_29  ( .a(\ne_42/AEQB [29]), .b(\ne_42/LTV [29]), .out(
        \ne_42/LTV2 [29]) );
  nand2 \ne_42/ULTI2_29  ( .a(\ne_42/LTV1 [29]), .b(\ne_42/LTV2 [29]), .out(
        \ne_42/LTV [30]) );
  xor2 \ne_42/UEQI_30  ( .a(final_floor_elevator2[30]), .b(requested_floor[30]), .out(n1783) );
  nand2 \ne_42/UGTI0_30  ( .a(n1782), .b(final_floor_elevator2[30]), .out(
        \ne_42/GTV1 [30]) );
  nand2 \ne_42/UGTI1_30  ( .a(\ne_42/AEQB [30]), .b(\ne_42/GTV [30]), .out(
        \ne_42/GTV2 [30]) );
  nand2 \ne_42/UGTI2_30  ( .a(\ne_42/GTV1 [30]), .b(\ne_42/GTV2 [30]), .out(
        \ne_42/GTV [31]) );
  nand2 \ne_42/ULTI0_30  ( .a(n1781), .b(requested_floor[30]), .out(
        \ne_42/LTV1 [30]) );
  nand2 \ne_42/ULTI1_30  ( .a(\ne_42/AEQB [30]), .b(\ne_42/LTV [30]), .out(
        \ne_42/LTV2 [30]) );
  nand2 \ne_42/ULTI2_30  ( .a(\ne_42/LTV1 [30]), .b(\ne_42/LTV2 [30]), .out(
        \ne_42/LTV [31]) );
  xor2 \ne_42/UEQI_31  ( .a(final_floor_elevator2[31]), .b(requested_floor[31]), .out(n1780) );
  nand2 \ne_42/UGTI0_31  ( .a(n1779), .b(final_floor_elevator2[31]), .out(
        \ne_42/GTV1 [31]) );
  nand2 \ne_42/UGTI1_31  ( .a(\ne_42/AEQB [31]), .b(\ne_42/GTV [31]), .out(
        \ne_42/GTV2 [31]) );
  nand2 \ne_42/UGTI2_31  ( .a(\ne_42/GTV1 [31]), .b(\ne_42/GTV2 [31]), .out(
        \ne_42/GTV [32]) );
  nand2 \ne_42/ULTI0_31  ( .a(n1778), .b(requested_floor[31]), .out(
        \ne_42/LTV1 [31]) );
  nand2 \ne_42/ULTI1_31  ( .a(\ne_42/AEQB [31]), .b(\ne_42/LTV [31]), .out(
        \ne_42/LTV2 [31]) );
  nand2 \ne_42/ULTI2_31  ( .a(\ne_42/LTV1 [31]), .b(\ne_42/LTV2 [31]), .out(
        \ne_42/LTV [32]) );
  xor2 \ne_42/UEQI_32  ( .a(final_floor_elevator2[32]), .b(requested_floor[32]), .out(n1777) );
  nand2 \ne_42/UGTI0_32  ( .a(n1776), .b(final_floor_elevator2[32]), .out(
        \ne_42/GTV1 [32]) );
  nand2 \ne_42/UGTI1_32  ( .a(\ne_42/AEQB [32]), .b(\ne_42/GTV [32]), .out(
        \ne_42/GTV2 [32]) );
  nand2 \ne_42/UGTI2_32  ( .a(\ne_42/GTV1 [32]), .b(\ne_42/GTV2 [32]), .out(
        \ne_42/GTV [33]) );
  nand2 \ne_42/ULTI0_32  ( .a(n1775), .b(requested_floor[32]), .out(
        \ne_42/LTV1 [32]) );
  nand2 \ne_42/ULTI1_32  ( .a(\ne_42/AEQB [32]), .b(\ne_42/LTV [32]), .out(
        \ne_42/LTV2 [32]) );
  nand2 \ne_42/ULTI2_32  ( .a(\ne_42/LTV1 [32]), .b(\ne_42/LTV2 [32]), .out(
        \ne_42/LTV [33]) );
  xor2 \ne_42/UEQI_33  ( .a(final_floor_elevator2[33]), .b(requested_floor[33]), .out(n1774) );
  nand2 \ne_42/UGTI0_33  ( .a(n1773), .b(final_floor_elevator2[33]), .out(
        \ne_42/GTV1 [33]) );
  nand2 \ne_42/UGTI1_33  ( .a(\ne_42/AEQB [33]), .b(\ne_42/GTV [33]), .out(
        \ne_42/GTV2 [33]) );
  nand2 \ne_42/UGTI2_33  ( .a(\ne_42/GTV1 [33]), .b(\ne_42/GTV2 [33]), .out(
        \ne_42/GTV [34]) );
  nand2 \ne_42/ULTI0_33  ( .a(n1772), .b(requested_floor[33]), .out(
        \ne_42/LTV1 [33]) );
  nand2 \ne_42/ULTI1_33  ( .a(\ne_42/AEQB [33]), .b(\ne_42/LTV [33]), .out(
        \ne_42/LTV2 [33]) );
  nand2 \ne_42/ULTI2_33  ( .a(\ne_42/LTV1 [33]), .b(\ne_42/LTV2 [33]), .out(
        \ne_42/LTV [34]) );
  xor2 \ne_42/UEQI_34  ( .a(final_floor_elevator2[34]), .b(requested_floor[34]), .out(n1771) );
  nand2 \ne_42/UGTI0_34  ( .a(n1770), .b(final_floor_elevator2[34]), .out(
        \ne_42/GTV1 [34]) );
  nand2 \ne_42/UGTI1_34  ( .a(\ne_42/AEQB [34]), .b(\ne_42/GTV [34]), .out(
        \ne_42/GTV2 [34]) );
  nand2 \ne_42/UGTI2_34  ( .a(\ne_42/GTV1 [34]), .b(\ne_42/GTV2 [34]), .out(
        \ne_42/GTV [35]) );
  nand2 \ne_42/ULTI0_34  ( .a(n1769), .b(requested_floor[34]), .out(
        \ne_42/LTV1 [34]) );
  nand2 \ne_42/ULTI1_34  ( .a(\ne_42/AEQB [34]), .b(\ne_42/LTV [34]), .out(
        \ne_42/LTV2 [34]) );
  nand2 \ne_42/ULTI2_34  ( .a(\ne_42/LTV1 [34]), .b(\ne_42/LTV2 [34]), .out(
        \ne_42/LTV [35]) );
  xor2 \ne_42/UEQI_35  ( .a(final_floor_elevator2[35]), .b(requested_floor[35]), .out(n1768) );
  nand2 \ne_42/UGTI0_35  ( .a(n1767), .b(final_floor_elevator2[35]), .out(
        \ne_42/GTV1 [35]) );
  nand2 \ne_42/UGTI1_35  ( .a(\ne_42/AEQB [35]), .b(\ne_42/GTV [35]), .out(
        \ne_42/GTV2 [35]) );
  nand2 \ne_42/UGTI2_35  ( .a(\ne_42/GTV1 [35]), .b(\ne_42/GTV2 [35]), .out(
        \ne_42/GTV [36]) );
  nand2 \ne_42/ULTI0_35  ( .a(n1766), .b(requested_floor[35]), .out(
        \ne_42/LTV1 [35]) );
  nand2 \ne_42/ULTI1_35  ( .a(\ne_42/AEQB [35]), .b(\ne_42/LTV [35]), .out(
        \ne_42/LTV2 [35]) );
  nand2 \ne_42/ULTI2_35  ( .a(\ne_42/LTV1 [35]), .b(\ne_42/LTV2 [35]), .out(
        \ne_42/LTV [36]) );
  xor2 \ne_42/UEQI_36  ( .a(final_floor_elevator2[36]), .b(requested_floor[36]), .out(n1765) );
  nand2 \ne_42/UGTI0_36  ( .a(n1764), .b(final_floor_elevator2[36]), .out(
        \ne_42/GTV1 [36]) );
  nand2 \ne_42/UGTI1_36  ( .a(\ne_42/AEQB [36]), .b(\ne_42/GTV [36]), .out(
        \ne_42/GTV2 [36]) );
  nand2 \ne_42/UGTI2_36  ( .a(\ne_42/GTV1 [36]), .b(\ne_42/GTV2 [36]), .out(
        \ne_42/GTV [37]) );
  nand2 \ne_42/ULTI0_36  ( .a(n1763), .b(requested_floor[36]), .out(
        \ne_42/LTV1 [36]) );
  nand2 \ne_42/ULTI1_36  ( .a(\ne_42/AEQB [36]), .b(\ne_42/LTV [36]), .out(
        \ne_42/LTV2 [36]) );
  nand2 \ne_42/ULTI2_36  ( .a(\ne_42/LTV1 [36]), .b(\ne_42/LTV2 [36]), .out(
        \ne_42/LTV [37]) );
  xor2 \ne_42/UEQI_37  ( .a(final_floor_elevator2[37]), .b(requested_floor[37]), .out(n1762) );
  nand2 \ne_42/UGTI0_37  ( .a(n1761), .b(final_floor_elevator2[37]), .out(
        \ne_42/GTV1 [37]) );
  nand2 \ne_42/UGTI1_37  ( .a(\ne_42/AEQB [37]), .b(\ne_42/GTV [37]), .out(
        \ne_42/GTV2 [37]) );
  nand2 \ne_42/UGTI2_37  ( .a(\ne_42/GTV1 [37]), .b(\ne_42/GTV2 [37]), .out(
        \ne_42/GTV [38]) );
  nand2 \ne_42/ULTI0_37  ( .a(n1760), .b(requested_floor[37]), .out(
        \ne_42/LTV1 [37]) );
  nand2 \ne_42/ULTI1_37  ( .a(\ne_42/AEQB [37]), .b(\ne_42/LTV [37]), .out(
        \ne_42/LTV2 [37]) );
  nand2 \ne_42/ULTI2_37  ( .a(\ne_42/LTV1 [37]), .b(\ne_42/LTV2 [37]), .out(
        \ne_42/LTV [38]) );
  xor2 \ne_42/UEQI_38  ( .a(final_floor_elevator2[38]), .b(requested_floor[38]), .out(n1759) );
  nand2 \ne_42/UGTI0_38  ( .a(n1758), .b(final_floor_elevator2[38]), .out(
        \ne_42/GTV1 [38]) );
  nand2 \ne_42/UGTI1_38  ( .a(\ne_42/AEQB [38]), .b(\ne_42/GTV [38]), .out(
        \ne_42/GTV2 [38]) );
  nand2 \ne_42/UGTI2_38  ( .a(\ne_42/GTV1 [38]), .b(\ne_42/GTV2 [38]), .out(
        \ne_42/GTV [39]) );
  nand2 \ne_42/ULTI0_38  ( .a(n1757), .b(requested_floor[38]), .out(
        \ne_42/LTV1 [38]) );
  nand2 \ne_42/ULTI1_38  ( .a(\ne_42/AEQB [38]), .b(\ne_42/LTV [38]), .out(
        \ne_42/LTV2 [38]) );
  nand2 \ne_42/ULTI2_38  ( .a(\ne_42/LTV1 [38]), .b(\ne_42/LTV2 [38]), .out(
        \ne_42/LTV [39]) );
  xor2 \ne_42/UEQI_39  ( .a(final_floor_elevator2[39]), .b(requested_floor[39]), .out(n1756) );
  nand2 \ne_42/UGTI0_39  ( .a(n1755), .b(final_floor_elevator2[39]), .out(
        \ne_42/GTV1 [39]) );
  nand2 \ne_42/UGTI1_39  ( .a(\ne_42/AEQB [39]), .b(\ne_42/GTV [39]), .out(
        \ne_42/GTV2 [39]) );
  nand2 \ne_42/UGTI2_39  ( .a(\ne_42/GTV1 [39]), .b(\ne_42/GTV2 [39]), .out(
        \ne_42/GTV [40]) );
  nand2 \ne_42/ULTI0_39  ( .a(n1754), .b(requested_floor[39]), .out(
        \ne_42/LTV1 [39]) );
  nand2 \ne_42/ULTI1_39  ( .a(\ne_42/AEQB [39]), .b(\ne_42/LTV [39]), .out(
        \ne_42/LTV2 [39]) );
  nand2 \ne_42/ULTI2_39  ( .a(\ne_42/LTV1 [39]), .b(\ne_42/LTV2 [39]), .out(
        \ne_42/LTV [40]) );
  xor2 \ne_42/UEQI_40  ( .a(final_floor_elevator2[40]), .b(requested_floor[40]), .out(n1753) );
  nand2 \ne_42/UGTI0_40  ( .a(n1752), .b(final_floor_elevator2[40]), .out(
        \ne_42/GTV1 [40]) );
  nand2 \ne_42/UGTI1_40  ( .a(\ne_42/AEQB [40]), .b(\ne_42/GTV [40]), .out(
        \ne_42/GTV2 [40]) );
  nand2 \ne_42/UGTI2_40  ( .a(\ne_42/GTV1 [40]), .b(\ne_42/GTV2 [40]), .out(
        \ne_42/GTV [41]) );
  nand2 \ne_42/ULTI0_40  ( .a(n1751), .b(requested_floor[40]), .out(
        \ne_42/LTV1 [40]) );
  nand2 \ne_42/ULTI1_40  ( .a(\ne_42/AEQB [40]), .b(\ne_42/LTV [40]), .out(
        \ne_42/LTV2 [40]) );
  nand2 \ne_42/ULTI2_40  ( .a(\ne_42/LTV1 [40]), .b(\ne_42/LTV2 [40]), .out(
        \ne_42/LTV [41]) );
  xor2 \ne_42/UEQI_41  ( .a(final_floor_elevator2[41]), .b(requested_floor[41]), .out(n1750) );
  nand2 \ne_42/UGTI0_41  ( .a(n1749), .b(final_floor_elevator2[41]), .out(
        \ne_42/GTV1 [41]) );
  nand2 \ne_42/UGTI1_41  ( .a(\ne_42/AEQB [41]), .b(\ne_42/GTV [41]), .out(
        \ne_42/GTV2 [41]) );
  nand2 \ne_42/UGTI2_41  ( .a(\ne_42/GTV1 [41]), .b(\ne_42/GTV2 [41]), .out(
        \ne_42/GTV [42]) );
  nand2 \ne_42/ULTI0_41  ( .a(n1748), .b(requested_floor[41]), .out(
        \ne_42/LTV1 [41]) );
  nand2 \ne_42/ULTI1_41  ( .a(\ne_42/AEQB [41]), .b(\ne_42/LTV [41]), .out(
        \ne_42/LTV2 [41]) );
  nand2 \ne_42/ULTI2_41  ( .a(\ne_42/LTV1 [41]), .b(\ne_42/LTV2 [41]), .out(
        \ne_42/LTV [42]) );
  xor2 \ne_42/UEQI_42  ( .a(final_floor_elevator2[42]), .b(requested_floor[42]), .out(n1747) );
  nand2 \ne_42/UGTI0_42  ( .a(n1746), .b(final_floor_elevator2[42]), .out(
        \ne_42/GTV1 [42]) );
  nand2 \ne_42/UGTI1_42  ( .a(\ne_42/AEQB [42]), .b(\ne_42/GTV [42]), .out(
        \ne_42/GTV2 [42]) );
  nand2 \ne_42/UGTI2_42  ( .a(\ne_42/GTV1 [42]), .b(\ne_42/GTV2 [42]), .out(
        \ne_42/GTV [43]) );
  nand2 \ne_42/ULTI0_42  ( .a(n1745), .b(requested_floor[42]), .out(
        \ne_42/LTV1 [42]) );
  nand2 \ne_42/ULTI1_42  ( .a(\ne_42/AEQB [42]), .b(\ne_42/LTV [42]), .out(
        \ne_42/LTV2 [42]) );
  nand2 \ne_42/ULTI2_42  ( .a(\ne_42/LTV1 [42]), .b(\ne_42/LTV2 [42]), .out(
        \ne_42/LTV [43]) );
  xor2 \ne_42/UEQI_43  ( .a(final_floor_elevator2[43]), .b(requested_floor[43]), .out(n1744) );
  nand2 \ne_42/UGTI0_43  ( .a(n1743), .b(final_floor_elevator2[43]), .out(
        \ne_42/GTV1 [43]) );
  nand2 \ne_42/UGTI1_43  ( .a(\ne_42/AEQB [43]), .b(\ne_42/GTV [43]), .out(
        \ne_42/GTV2 [43]) );
  nand2 \ne_42/UGTI2_43  ( .a(\ne_42/GTV1 [43]), .b(\ne_42/GTV2 [43]), .out(
        \ne_42/GTV [44]) );
  nand2 \ne_42/ULTI0_43  ( .a(n1742), .b(requested_floor[43]), .out(
        \ne_42/LTV1 [43]) );
  nand2 \ne_42/ULTI1_43  ( .a(\ne_42/AEQB [43]), .b(\ne_42/LTV [43]), .out(
        \ne_42/LTV2 [43]) );
  nand2 \ne_42/ULTI2_43  ( .a(\ne_42/LTV1 [43]), .b(\ne_42/LTV2 [43]), .out(
        \ne_42/LTV [44]) );
  xor2 \ne_42/UEQI_44  ( .a(final_floor_elevator2[44]), .b(requested_floor[44]), .out(n1741) );
  nand2 \ne_42/UGTI0_44  ( .a(n1740), .b(final_floor_elevator2[44]), .out(
        \ne_42/GTV1 [44]) );
  nand2 \ne_42/UGTI1_44  ( .a(\ne_42/AEQB [44]), .b(\ne_42/GTV [44]), .out(
        \ne_42/GTV2 [44]) );
  nand2 \ne_42/UGTI2_44  ( .a(\ne_42/GTV1 [44]), .b(\ne_42/GTV2 [44]), .out(
        \ne_42/GTV [45]) );
  nand2 \ne_42/ULTI0_44  ( .a(n1739), .b(requested_floor[44]), .out(
        \ne_42/LTV1 [44]) );
  nand2 \ne_42/ULTI1_44  ( .a(\ne_42/AEQB [44]), .b(\ne_42/LTV [44]), .out(
        \ne_42/LTV2 [44]) );
  nand2 \ne_42/ULTI2_44  ( .a(\ne_42/LTV1 [44]), .b(\ne_42/LTV2 [44]), .out(
        \ne_42/LTV [45]) );
  xor2 \ne_42/UEQI_45  ( .a(final_floor_elevator2[45]), .b(requested_floor[45]), .out(n1738) );
  nand2 \ne_42/UGTI0_45  ( .a(n1737), .b(final_floor_elevator2[45]), .out(
        \ne_42/GTV1 [45]) );
  nand2 \ne_42/UGTI1_45  ( .a(\ne_42/AEQB [45]), .b(\ne_42/GTV [45]), .out(
        \ne_42/GTV2 [45]) );
  nand2 \ne_42/UGTI2_45  ( .a(\ne_42/GTV1 [45]), .b(\ne_42/GTV2 [45]), .out(
        \ne_42/GTV [46]) );
  nand2 \ne_42/ULTI0_45  ( .a(n1736), .b(requested_floor[45]), .out(
        \ne_42/LTV1 [45]) );
  nand2 \ne_42/ULTI1_45  ( .a(\ne_42/AEQB [45]), .b(\ne_42/LTV [45]), .out(
        \ne_42/LTV2 [45]) );
  nand2 \ne_42/ULTI2_45  ( .a(\ne_42/LTV1 [45]), .b(\ne_42/LTV2 [45]), .out(
        \ne_42/LTV [46]) );
  xor2 \ne_42/UEQI_46  ( .a(final_floor_elevator2[46]), .b(requested_floor[46]), .out(n1735) );
  nand2 \ne_42/UGTI0_46  ( .a(n1734), .b(final_floor_elevator2[46]), .out(
        \ne_42/GTV1 [46]) );
  nand2 \ne_42/UGTI1_46  ( .a(\ne_42/AEQB [46]), .b(\ne_42/GTV [46]), .out(
        \ne_42/GTV2 [46]) );
  nand2 \ne_42/UGTI2_46  ( .a(\ne_42/GTV1 [46]), .b(\ne_42/GTV2 [46]), .out(
        \ne_42/GTV [47]) );
  nand2 \ne_42/ULTI0_46  ( .a(n1733), .b(requested_floor[46]), .out(
        \ne_42/LTV1 [46]) );
  nand2 \ne_42/ULTI1_46  ( .a(\ne_42/AEQB [46]), .b(\ne_42/LTV [46]), .out(
        \ne_42/LTV2 [46]) );
  nand2 \ne_42/ULTI2_46  ( .a(\ne_42/LTV1 [46]), .b(\ne_42/LTV2 [46]), .out(
        \ne_42/LTV [47]) );
  xor2 \ne_42/UEQI_47  ( .a(final_floor_elevator2[47]), .b(requested_floor[47]), .out(n1732) );
  nand2 \ne_42/UGTI0_47  ( .a(n1731), .b(final_floor_elevator2[47]), .out(
        \ne_42/GTV1 [47]) );
  nand2 \ne_42/UGTI1_47  ( .a(\ne_42/AEQB [47]), .b(\ne_42/GTV [47]), .out(
        \ne_42/GTV2 [47]) );
  nand2 \ne_42/UGTI2_47  ( .a(\ne_42/GTV1 [47]), .b(\ne_42/GTV2 [47]), .out(
        \ne_42/GTV [48]) );
  nand2 \ne_42/ULTI0_47  ( .a(n1730), .b(requested_floor[47]), .out(
        \ne_42/LTV1 [47]) );
  nand2 \ne_42/ULTI1_47  ( .a(\ne_42/AEQB [47]), .b(\ne_42/LTV [47]), .out(
        \ne_42/LTV2 [47]) );
  nand2 \ne_42/ULTI2_47  ( .a(\ne_42/LTV1 [47]), .b(\ne_42/LTV2 [47]), .out(
        \ne_42/LTV [48]) );
  xor2 \ne_42/UEQI_48  ( .a(final_floor_elevator2[48]), .b(requested_floor[48]), .out(n1729) );
  nand2 \ne_42/UGTI0_48  ( .a(n1728), .b(final_floor_elevator2[48]), .out(
        \ne_42/GTV1 [48]) );
  nand2 \ne_42/UGTI1_48  ( .a(\ne_42/AEQB [48]), .b(\ne_42/GTV [48]), .out(
        \ne_42/GTV2 [48]) );
  nand2 \ne_42/UGTI2_48  ( .a(\ne_42/GTV1 [48]), .b(\ne_42/GTV2 [48]), .out(
        \ne_42/GTV [49]) );
  nand2 \ne_42/ULTI0_48  ( .a(n1727), .b(requested_floor[48]), .out(
        \ne_42/LTV1 [48]) );
  nand2 \ne_42/ULTI1_48  ( .a(\ne_42/AEQB [48]), .b(\ne_42/LTV [48]), .out(
        \ne_42/LTV2 [48]) );
  nand2 \ne_42/ULTI2_48  ( .a(\ne_42/LTV1 [48]), .b(\ne_42/LTV2 [48]), .out(
        \ne_42/LTV [49]) );
  xor2 \ne_42/UEQI_49  ( .a(final_floor_elevator2[49]), .b(requested_floor[49]), .out(n1726) );
  nand2 \ne_42/UGTI0_49  ( .a(n1725), .b(final_floor_elevator2[49]), .out(
        \ne_42/GTV1 [49]) );
  nand2 \ne_42/UGTI1_49  ( .a(\ne_42/AEQB [49]), .b(\ne_42/GTV [49]), .out(
        \ne_42/GTV2 [49]) );
  nand2 \ne_42/UGTI2_49  ( .a(\ne_42/GTV1 [49]), .b(\ne_42/GTV2 [49]), .out(
        \ne_42/GTV [50]) );
  nand2 \ne_42/ULTI0_49  ( .a(n1724), .b(requested_floor[49]), .out(
        \ne_42/LTV1 [49]) );
  nand2 \ne_42/ULTI1_49  ( .a(\ne_42/AEQB [49]), .b(\ne_42/LTV [49]), .out(
        \ne_42/LTV2 [49]) );
  nand2 \ne_42/ULTI2_49  ( .a(\ne_42/LTV1 [49]), .b(\ne_42/LTV2 [49]), .out(
        \ne_42/LTV [50]) );
  xor2 \ne_42/UEQI_50  ( .a(final_floor_elevator2[50]), .b(requested_floor[50]), .out(n1723) );
  nand2 \ne_42/UGTI0_50  ( .a(n1722), .b(final_floor_elevator2[50]), .out(
        \ne_42/GTV1 [50]) );
  nand2 \ne_42/UGTI1_50  ( .a(\ne_42/AEQB [50]), .b(\ne_42/GTV [50]), .out(
        \ne_42/GTV2 [50]) );
  nand2 \ne_42/UGTI2_50  ( .a(\ne_42/GTV1 [50]), .b(\ne_42/GTV2 [50]), .out(
        \ne_42/GTV [51]) );
  nand2 \ne_42/ULTI0_50  ( .a(n1721), .b(requested_floor[50]), .out(
        \ne_42/LTV1 [50]) );
  nand2 \ne_42/ULTI1_50  ( .a(\ne_42/AEQB [50]), .b(\ne_42/LTV [50]), .out(
        \ne_42/LTV2 [50]) );
  nand2 \ne_42/ULTI2_50  ( .a(\ne_42/LTV1 [50]), .b(\ne_42/LTV2 [50]), .out(
        \ne_42/LTV [51]) );
  xor2 \ne_42/UEQI_51  ( .a(final_floor_elevator2[51]), .b(requested_floor[51]), .out(n1720) );
  nand2 \ne_42/UGTI0_51  ( .a(n1719), .b(final_floor_elevator2[51]), .out(
        \ne_42/GTV1 [51]) );
  nand2 \ne_42/UGTI1_51  ( .a(\ne_42/AEQB [51]), .b(\ne_42/GTV [51]), .out(
        \ne_42/GTV2 [51]) );
  nand2 \ne_42/UGTI2_51  ( .a(\ne_42/GTV1 [51]), .b(\ne_42/GTV2 [51]), .out(
        \ne_42/GTV [52]) );
  nand2 \ne_42/ULTI0_51  ( .a(n1718), .b(requested_floor[51]), .out(
        \ne_42/LTV1 [51]) );
  nand2 \ne_42/ULTI1_51  ( .a(\ne_42/AEQB [51]), .b(\ne_42/LTV [51]), .out(
        \ne_42/LTV2 [51]) );
  nand2 \ne_42/ULTI2_51  ( .a(\ne_42/LTV1 [51]), .b(\ne_42/LTV2 [51]), .out(
        \ne_42/LTV [52]) );
  xor2 \ne_42/UEQI_52  ( .a(final_floor_elevator2[52]), .b(requested_floor[52]), .out(n1717) );
  nand2 \ne_42/UGTI0_52  ( .a(n1716), .b(final_floor_elevator2[52]), .out(
        \ne_42/GTV1 [52]) );
  nand2 \ne_42/UGTI1_52  ( .a(\ne_42/AEQB [52]), .b(\ne_42/GTV [52]), .out(
        \ne_42/GTV2 [52]) );
  nand2 \ne_42/UGTI2_52  ( .a(\ne_42/GTV1 [52]), .b(\ne_42/GTV2 [52]), .out(
        \ne_42/GTV [53]) );
  nand2 \ne_42/ULTI0_52  ( .a(n1715), .b(requested_floor[52]), .out(
        \ne_42/LTV1 [52]) );
  nand2 \ne_42/ULTI1_52  ( .a(\ne_42/AEQB [52]), .b(\ne_42/LTV [52]), .out(
        \ne_42/LTV2 [52]) );
  nand2 \ne_42/ULTI2_52  ( .a(\ne_42/LTV1 [52]), .b(\ne_42/LTV2 [52]), .out(
        \ne_42/LTV [53]) );
  xor2 \ne_42/UEQI_53  ( .a(final_floor_elevator2[53]), .b(requested_floor[53]), .out(n1714) );
  nand2 \ne_42/UGTI0_53  ( .a(n1713), .b(final_floor_elevator2[53]), .out(
        \ne_42/GTV1 [53]) );
  nand2 \ne_42/UGTI1_53  ( .a(\ne_42/AEQB [53]), .b(\ne_42/GTV [53]), .out(
        \ne_42/GTV2 [53]) );
  nand2 \ne_42/UGTI2_53  ( .a(\ne_42/GTV1 [53]), .b(\ne_42/GTV2 [53]), .out(
        \ne_42/GTV [54]) );
  nand2 \ne_42/ULTI0_53  ( .a(n1712), .b(requested_floor[53]), .out(
        \ne_42/LTV1 [53]) );
  nand2 \ne_42/ULTI1_53  ( .a(\ne_42/AEQB [53]), .b(\ne_42/LTV [53]), .out(
        \ne_42/LTV2 [53]) );
  nand2 \ne_42/ULTI2_53  ( .a(\ne_42/LTV1 [53]), .b(\ne_42/LTV2 [53]), .out(
        \ne_42/LTV [54]) );
  xor2 \ne_42/UEQI_54  ( .a(final_floor_elevator2[54]), .b(requested_floor[54]), .out(n1711) );
  nand2 \ne_42/UGTI0_54  ( .a(n1710), .b(final_floor_elevator2[54]), .out(
        \ne_42/GTV1 [54]) );
  nand2 \ne_42/UGTI1_54  ( .a(\ne_42/AEQB [54]), .b(\ne_42/GTV [54]), .out(
        \ne_42/GTV2 [54]) );
  nand2 \ne_42/UGTI2_54  ( .a(\ne_42/GTV1 [54]), .b(\ne_42/GTV2 [54]), .out(
        \ne_42/GTV [55]) );
  nand2 \ne_42/ULTI0_54  ( .a(n1709), .b(requested_floor[54]), .out(
        \ne_42/LTV1 [54]) );
  nand2 \ne_42/ULTI1_54  ( .a(\ne_42/AEQB [54]), .b(\ne_42/LTV [54]), .out(
        \ne_42/LTV2 [54]) );
  nand2 \ne_42/ULTI2_54  ( .a(\ne_42/LTV1 [54]), .b(\ne_42/LTV2 [54]), .out(
        \ne_42/LTV [55]) );
  xor2 \ne_42/UEQI_55  ( .a(final_floor_elevator2[55]), .b(requested_floor[55]), .out(n1708) );
  nand2 \ne_42/UGTI0_55  ( .a(n1707), .b(final_floor_elevator2[55]), .out(
        \ne_42/GTV1 [55]) );
  nand2 \ne_42/UGTI1_55  ( .a(\ne_42/AEQB [55]), .b(\ne_42/GTV [55]), .out(
        \ne_42/GTV2 [55]) );
  nand2 \ne_42/UGTI2_55  ( .a(\ne_42/GTV1 [55]), .b(\ne_42/GTV2 [55]), .out(
        \ne_42/GTV [56]) );
  nand2 \ne_42/ULTI0_55  ( .a(n1706), .b(requested_floor[55]), .out(
        \ne_42/LTV1 [55]) );
  nand2 \ne_42/ULTI1_55  ( .a(\ne_42/AEQB [55]), .b(\ne_42/LTV [55]), .out(
        \ne_42/LTV2 [55]) );
  nand2 \ne_42/ULTI2_55  ( .a(\ne_42/LTV1 [55]), .b(\ne_42/LTV2 [55]), .out(
        \ne_42/LTV [56]) );
  xor2 \ne_42/UEQI_56  ( .a(final_floor_elevator2[56]), .b(requested_floor[56]), .out(n1705) );
  nand2 \ne_42/UGTI0_56  ( .a(n1704), .b(final_floor_elevator2[56]), .out(
        \ne_42/GTV1 [56]) );
  nand2 \ne_42/UGTI1_56  ( .a(\ne_42/AEQB [56]), .b(\ne_42/GTV [56]), .out(
        \ne_42/GTV2 [56]) );
  nand2 \ne_42/UGTI2_56  ( .a(\ne_42/GTV1 [56]), .b(\ne_42/GTV2 [56]), .out(
        \ne_42/GTV [57]) );
  nand2 \ne_42/ULTI0_56  ( .a(n1703), .b(requested_floor[56]), .out(
        \ne_42/LTV1 [56]) );
  nand2 \ne_42/ULTI1_56  ( .a(\ne_42/AEQB [56]), .b(\ne_42/LTV [56]), .out(
        \ne_42/LTV2 [56]) );
  nand2 \ne_42/ULTI2_56  ( .a(\ne_42/LTV1 [56]), .b(\ne_42/LTV2 [56]), .out(
        \ne_42/LTV [57]) );
  xor2 \ne_42/UEQI_57  ( .a(final_floor_elevator2[57]), .b(requested_floor[57]), .out(n1702) );
  nand2 \ne_42/UGTI0_57  ( .a(n1701), .b(final_floor_elevator2[57]), .out(
        \ne_42/GTV1 [57]) );
  nand2 \ne_42/UGTI1_57  ( .a(\ne_42/AEQB [57]), .b(\ne_42/GTV [57]), .out(
        \ne_42/GTV2 [57]) );
  nand2 \ne_42/UGTI2_57  ( .a(\ne_42/GTV1 [57]), .b(\ne_42/GTV2 [57]), .out(
        \ne_42/GTV [58]) );
  nand2 \ne_42/ULTI0_57  ( .a(n1700), .b(requested_floor[57]), .out(
        \ne_42/LTV1 [57]) );
  nand2 \ne_42/ULTI1_57  ( .a(\ne_42/AEQB [57]), .b(\ne_42/LTV [57]), .out(
        \ne_42/LTV2 [57]) );
  nand2 \ne_42/ULTI2_57  ( .a(\ne_42/LTV1 [57]), .b(\ne_42/LTV2 [57]), .out(
        \ne_42/LTV [58]) );
  xor2 \ne_42/UEQI_58  ( .a(final_floor_elevator2[58]), .b(requested_floor[58]), .out(n1699) );
  nand2 \ne_42/UGTI0_58  ( .a(n1698), .b(final_floor_elevator2[58]), .out(
        \ne_42/GTV1 [58]) );
  nand2 \ne_42/UGTI1_58  ( .a(\ne_42/AEQB [58]), .b(\ne_42/GTV [58]), .out(
        \ne_42/GTV2 [58]) );
  nand2 \ne_42/UGTI2_58  ( .a(\ne_42/GTV1 [58]), .b(\ne_42/GTV2 [58]), .out(
        \ne_42/GTV [59]) );
  nand2 \ne_42/ULTI0_58  ( .a(n1697), .b(requested_floor[58]), .out(
        \ne_42/LTV1 [58]) );
  nand2 \ne_42/ULTI1_58  ( .a(\ne_42/AEQB [58]), .b(\ne_42/LTV [58]), .out(
        \ne_42/LTV2 [58]) );
  nand2 \ne_42/ULTI2_58  ( .a(\ne_42/LTV1 [58]), .b(\ne_42/LTV2 [58]), .out(
        \ne_42/LTV [59]) );
  xor2 \ne_42/UEQI_59  ( .a(final_floor_elevator2[59]), .b(requested_floor[59]), .out(n1696) );
  nand2 \ne_42/UGTI0_59  ( .a(n1695), .b(final_floor_elevator2[59]), .out(
        \ne_42/GTV1 [59]) );
  nand2 \ne_42/UGTI1_59  ( .a(\ne_42/AEQB [59]), .b(\ne_42/GTV [59]), .out(
        \ne_42/GTV2 [59]) );
  nand2 \ne_42/UGTI2_59  ( .a(\ne_42/GTV1 [59]), .b(\ne_42/GTV2 [59]), .out(
        \ne_42/GTV [60]) );
  nand2 \ne_42/ULTI0_59  ( .a(n1694), .b(requested_floor[59]), .out(
        \ne_42/LTV1 [59]) );
  nand2 \ne_42/ULTI1_59  ( .a(\ne_42/AEQB [59]), .b(\ne_42/LTV [59]), .out(
        \ne_42/LTV2 [59]) );
  nand2 \ne_42/ULTI2_59  ( .a(\ne_42/LTV1 [59]), .b(\ne_42/LTV2 [59]), .out(
        \ne_42/LTV [60]) );
  xor2 \ne_42/UEQI_60  ( .a(final_floor_elevator2[60]), .b(requested_floor[60]), .out(n1693) );
  nand2 \ne_42/UGTI0_60  ( .a(n1692), .b(final_floor_elevator2[60]), .out(
        \ne_42/GTV1 [60]) );
  nand2 \ne_42/UGTI1_60  ( .a(\ne_42/AEQB [60]), .b(\ne_42/GTV [60]), .out(
        \ne_42/GTV2 [60]) );
  nand2 \ne_42/UGTI2_60  ( .a(\ne_42/GTV1 [60]), .b(\ne_42/GTV2 [60]), .out(
        \ne_42/GTV [61]) );
  nand2 \ne_42/ULTI0_60  ( .a(n1691), .b(requested_floor[60]), .out(
        \ne_42/LTV1 [60]) );
  nand2 \ne_42/ULTI1_60  ( .a(\ne_42/AEQB [60]), .b(\ne_42/LTV [60]), .out(
        \ne_42/LTV2 [60]) );
  nand2 \ne_42/ULTI2_60  ( .a(\ne_42/LTV1 [60]), .b(\ne_42/LTV2 [60]), .out(
        \ne_42/LTV [61]) );
  xor2 \ne_42/UEQI_61  ( .a(final_floor_elevator2[61]), .b(requested_floor[61]), .out(n1690) );
  nand2 \ne_42/UGTI0_61  ( .a(n1689), .b(final_floor_elevator2[61]), .out(
        \ne_42/GTV1 [61]) );
  nand2 \ne_42/UGTI1_61  ( .a(\ne_42/AEQB [61]), .b(\ne_42/GTV [61]), .out(
        \ne_42/GTV2 [61]) );
  nand2 \ne_42/UGTI2_61  ( .a(\ne_42/GTV1 [61]), .b(\ne_42/GTV2 [61]), .out(
        \ne_42/GTV [62]) );
  nand2 \ne_42/ULTI0_61  ( .a(n1688), .b(requested_floor[61]), .out(
        \ne_42/LTV1 [61]) );
  nand2 \ne_42/ULTI1_61  ( .a(\ne_42/AEQB [61]), .b(\ne_42/LTV [61]), .out(
        \ne_42/LTV2 [61]) );
  nand2 \ne_42/ULTI2_61  ( .a(\ne_42/LTV1 [61]), .b(\ne_42/LTV2 [61]), .out(
        \ne_42/LTV [62]) );
  xor2 \ne_42/UEQI_62  ( .a(final_floor_elevator2[62]), .b(requested_floor[62]), .out(n1687) );
  nand2 \ne_42/UGTI0_62  ( .a(n1686), .b(final_floor_elevator2[62]), .out(
        \ne_42/GTV1 [62]) );
  nand2 \ne_42/UGTI1_62  ( .a(\ne_42/AEQB [62]), .b(\ne_42/GTV [62]), .out(
        \ne_42/GTV2 [62]) );
  nand2 \ne_42/UGTI2_62  ( .a(\ne_42/GTV1 [62]), .b(\ne_42/GTV2 [62]), .out(
        \ne_42/GTV [63]) );
  nand2 \ne_42/ULTI0_62  ( .a(n1685), .b(requested_floor[62]), .out(
        \ne_42/LTV1 [62]) );
  nand2 \ne_42/ULTI1_62  ( .a(\ne_42/AEQB [62]), .b(\ne_42/LTV [62]), .out(
        \ne_42/LTV2 [62]) );
  nand2 \ne_42/ULTI2_62  ( .a(\ne_42/LTV1 [62]), .b(\ne_42/LTV2 [62]), .out(
        \ne_42/LTV [63]) );
  inv U1169 ( .in(n1493), .out(n1431) );
  inv U1170 ( .in(n1493), .out(n1432) );
  inv U1171 ( .in(n1492), .out(n1433) );
  inv U1172 ( .in(n1492), .out(n1434) );
  inv U1173 ( .in(n1492), .out(n1435) );
  inv U1174 ( .in(n1491), .out(n1436) );
  inv U1175 ( .in(n1491), .out(n1437) );
  inv U1176 ( .in(n1491), .out(n1438) );
  inv U1177 ( .in(n1490), .out(n1439) );
  inv U1178 ( .in(n1490), .out(n1440) );
  inv U1179 ( .in(n1490), .out(n1441) );
  inv U1180 ( .in(n1489), .out(n1442) );
  inv U1181 ( .in(n1489), .out(n1443) );
  inv U1182 ( .in(n1489), .out(n1444) );
  inv U1183 ( .in(n1488), .out(n1445) );
  inv U1184 ( .in(n1488), .out(n1446) );
  inv U1185 ( .in(n1488), .out(n1447) );
  inv U1186 ( .in(n1487), .out(n1448) );
  inv U1187 ( .in(n1487), .out(n1449) );
  inv U1188 ( .in(n1487), .out(n1450) );
  inv U1189 ( .in(n1486), .out(n1451) );
  inv U1190 ( .in(n1486), .out(n1452) );
  inv U1191 ( .in(n1486), .out(n1453) );
  inv U1192 ( .in(n1485), .out(n1454) );
  inv U1193 ( .in(n1485), .out(n1455) );
  inv U1194 ( .in(n1485), .out(n1456) );
  inv U1195 ( .in(n1484), .out(n1457) );
  inv U1196 ( .in(n1484), .out(n1458) );
  inv U1197 ( .in(n1484), .out(n1459) );
  inv U1198 ( .in(n1483), .out(n1460) );
  inv U1199 ( .in(n1483), .out(n1461) );
  inv U1200 ( .in(n1483), .out(n1462) );
  inv U1201 ( .in(n1482), .out(n1463) );
  inv U1202 ( .in(n1482), .out(n1464) );
  inv U1203 ( .in(n1482), .out(n1465) );
  inv U1204 ( .in(n1481), .out(n1466) );
  inv U1205 ( .in(n1481), .out(n1467) );
  inv U1206 ( .in(n1481), .out(n1468) );
  inv U1207 ( .in(n1480), .out(n1469) );
  inv U1208 ( .in(n1480), .out(n1470) );
  inv U1209 ( .in(n1480), .out(n1471) );
  inv U1210 ( .in(n1479), .out(n1472) );
  inv U1211 ( .in(n1479), .out(n1473) );
  inv U1212 ( .in(n1479), .out(n1474) );
  inv U1213 ( .in(n1478), .out(n1475) );
  inv U1214 ( .in(n1478), .out(n1476) );
  inv U1215 ( .in(n1478), .out(n1477) );
  inv U1216 ( .in(n1499), .out(n1478) );
  inv U1217 ( .in(n1498), .out(n1479) );
  inv U1218 ( .in(n1498), .out(n1480) );
  inv U1219 ( .in(n1498), .out(n1481) );
  inv U1220 ( .in(n1497), .out(n1482) );
  inv U1221 ( .in(n1497), .out(n1483) );
  inv U1222 ( .in(n1497), .out(n1484) );
  inv U1223 ( .in(n1496), .out(n1485) );
  inv U1224 ( .in(n1496), .out(n1486) );
  inv U1225 ( .in(n1496), .out(n1487) );
  inv U1226 ( .in(n1495), .out(n1488) );
  inv U1227 ( .in(n1495), .out(n1489) );
  inv U1228 ( .in(n1495), .out(n1490) );
  inv U1229 ( .in(n1494), .out(n1491) );
  inv U1230 ( .in(n1494), .out(n1492) );
  inv U1231 ( .in(n1494), .out(n1493) );
  inv U1232 ( .in(n1501), .out(n1494) );
  inv U1233 ( .in(n1501), .out(n1495) );
  inv U1234 ( .in(n1501), .out(n1496) );
  inv U1235 ( .in(n1500), .out(n1497) );
  inv U1236 ( .in(n1500), .out(n1498) );
  inv U1237 ( .in(n1500), .out(n1499) );
  inv U1238 ( .in(N360), .out(n1500) );
  inv U1239 ( .in(N360), .out(n1501) );
  inv U1240 ( .in(n1473), .out(n1502) );
  inv U1241 ( .in(n1474), .out(n1503) );
  inv U1242 ( .in(n1474), .out(n1504) );
  inv U1243 ( .in(n1474), .out(n1505) );
  inv U1244 ( .in(n1475), .out(n1506) );
  inv U1245 ( .in(n1475), .out(n1507) );
  inv U1246 ( .in(n1475), .out(n1508) );
  inv U1247 ( .in(n1476), .out(n1509) );
  inv U1248 ( .in(n1476), .out(n1510) );
  inv U1249 ( .in(n1476), .out(n1511) );
  inv U1250 ( .in(n1477), .out(n1512) );
  inv U1251 ( .in(n1575), .out(n1513) );
  inv U1252 ( .in(n1575), .out(n1514) );
  inv U1253 ( .in(n1574), .out(n1515) );
  inv U1254 ( .in(n1574), .out(n1516) );
  inv U1255 ( .in(n1574), .out(n1517) );
  inv U1256 ( .in(n1573), .out(n1518) );
  inv U1257 ( .in(n1573), .out(n1519) );
  inv U1258 ( .in(n1573), .out(n1520) );
  inv U1259 ( .in(n1572), .out(n1521) );
  inv U1260 ( .in(n1572), .out(n1522) );
  inv U1261 ( .in(n1572), .out(n1523) );
  inv U1262 ( .in(n1571), .out(n1524) );
  inv U1263 ( .in(n1571), .out(n1525) );
  inv U1264 ( .in(n1571), .out(n1526) );
  inv U1265 ( .in(n1570), .out(n1527) );
  inv U1266 ( .in(n1570), .out(n1528) );
  inv U1267 ( .in(n1570), .out(n1529) );
  inv U1268 ( .in(n1569), .out(n1530) );
  inv U1269 ( .in(n1569), .out(n1531) );
  inv U1270 ( .in(n1569), .out(n1532) );
  inv U1271 ( .in(n1568), .out(n1533) );
  inv U1272 ( .in(n1568), .out(n1534) );
  inv U1273 ( .in(n1568), .out(n1535) );
  inv U1274 ( .in(n1567), .out(n1536) );
  inv U1275 ( .in(n1567), .out(n1537) );
  inv U1276 ( .in(n1567), .out(n1538) );
  inv U1277 ( .in(n1566), .out(n1539) );
  inv U1278 ( .in(n1566), .out(n1540) );
  inv U1279 ( .in(n1566), .out(n1541) );
  inv U1280 ( .in(n1565), .out(n1542) );
  inv U1281 ( .in(n1565), .out(n1543) );
  inv U1282 ( .in(n1565), .out(n1544) );
  inv U1283 ( .in(n1564), .out(n1545) );
  inv U1284 ( .in(n1564), .out(n1546) );
  inv U1285 ( .in(n1564), .out(n1547) );
  inv U1286 ( .in(n1563), .out(n1548) );
  inv U1287 ( .in(n1563), .out(n1549) );
  inv U1288 ( .in(n1563), .out(n1550) );
  inv U1289 ( .in(n1562), .out(n1551) );
  inv U1290 ( .in(n1562), .out(n1552) );
  inv U1291 ( .in(n1562), .out(n1553) );
  inv U1292 ( .in(n1561), .out(n1554) );
  inv U1293 ( .in(n1561), .out(n1555) );
  inv U1294 ( .in(n1561), .out(n1556) );
  inv U1295 ( .in(n1560), .out(n1557) );
  inv U1296 ( .in(n1560), .out(n1558) );
  inv U1297 ( .in(n1560), .out(n1559) );
  inv U1298 ( .in(n1581), .out(n1560) );
  inv U1299 ( .in(n1580), .out(n1561) );
  inv U1300 ( .in(n1580), .out(n1562) );
  inv U1301 ( .in(n1580), .out(n1563) );
  inv U1302 ( .in(n1579), .out(n1564) );
  inv U1303 ( .in(n1579), .out(n1565) );
  inv U1304 ( .in(n1579), .out(n1566) );
  inv U1305 ( .in(n1578), .out(n1567) );
  inv U1306 ( .in(n1578), .out(n1568) );
  inv U1307 ( .in(n1578), .out(n1569) );
  inv U1308 ( .in(n1577), .out(n1570) );
  inv U1309 ( .in(n1577), .out(n1571) );
  inv U1310 ( .in(n1577), .out(n1572) );
  inv U1311 ( .in(n1576), .out(n1573) );
  inv U1312 ( .in(n1576), .out(n1574) );
  inv U1313 ( .in(n1576), .out(n1575) );
  inv U1314 ( .in(n1583), .out(n1576) );
  inv U1315 ( .in(n1583), .out(n1577) );
  inv U1316 ( .in(n1583), .out(n1578) );
  inv U1317 ( .in(n1582), .out(n1579) );
  inv U1318 ( .in(n1582), .out(n1580) );
  inv U1319 ( .in(n1582), .out(n1581) );
  inv U1320 ( .in(N76), .out(n1582) );
  inv U1321 ( .in(N76), .out(n1583) );
  inv U1322 ( .in(n1555), .out(n1584) );
  inv U1323 ( .in(n1556), .out(n1585) );
  inv U1324 ( .in(n1556), .out(n1586) );
  inv U1325 ( .in(n1556), .out(n1587) );
  inv U1326 ( .in(n1557), .out(n1588) );
  inv U1327 ( .in(n1557), .out(n1589) );
  inv U1328 ( .in(n1557), .out(n1590) );
  inv U1329 ( .in(n1558), .out(n1591) );
  inv U1330 ( .in(n1558), .out(n1592) );
  inv U1331 ( .in(n1558), .out(n1593) );
  inv U1332 ( .in(n1559), .out(n1594) );
  inv U1333 ( .in(n1617), .out(n1595) );
  inv U1334 ( .in(n1617), .out(n1596) );
  inv U1335 ( .in(n1616), .out(n1597) );
  inv U1336 ( .in(n1616), .out(n1598) );
  inv U1337 ( .in(n1616), .out(n1599) );
  inv U1338 ( .in(n1615), .out(n1600) );
  inv U1339 ( .in(n1615), .out(n1601) );
  inv U1340 ( .in(n1615), .out(n1602) );
  inv U1341 ( .in(n1614), .out(n1603) );
  inv U1342 ( .in(n1614), .out(n1604) );
  inv U1343 ( .in(n1614), .out(n1605) );
  inv U1344 ( .in(n1613), .out(n1606) );
  inv U1345 ( .in(n1613), .out(n1607) );
  inv U1346 ( .in(n1613), .out(n1608) );
  inv U1347 ( .in(n1612), .out(n1609) );
  inv U1348 ( .in(n1612), .out(n1610) );
  inv U1349 ( .in(n1612), .out(n1611) );
  inv U1350 ( .in(reset_elevator2), .out(n1612) );
  inv U1351 ( .in(reset_elevator2), .out(n1613) );
  inv U1352 ( .in(reset_elevator2), .out(n1614) );
  inv U1353 ( .in(reset_elevator2), .out(n1615) );
  inv U1354 ( .in(reset_elevator2), .out(n1616) );
  inv U1355 ( .in(reset_elevator2), .out(n1617) );
  inv U1356 ( .in(reset_elevator2), .out(n1618) );
  inv U1357 ( .in(reset_elevator2), .out(n1619) );
  inv U1358 ( .in(reset_elevator2), .out(n1620) );
  inv U1359 ( .in(reset_elevator2), .out(n1621) );
  inv U1360 ( .in(reset_elevator2), .out(n1622) );
  inv U1361 ( .in(reset_elevator2), .out(n1623) );
  inv U1362 ( .in(reset_elevator2), .out(n1624) );
  inv U1363 ( .in(reset_elevator2), .out(n1625) );
  inv U1364 ( .in(reset_elevator2), .out(n1626) );
  inv U1365 ( .in(reset_elevator2), .out(n1627) );
  inv U1366 ( .in(reset_elevator2), .out(n1628) );
  inv U1367 ( .in(reset_elevator2), .out(n1629) );
  inv U1368 ( .in(reset_elevator2), .out(n1630) );
  inv U1369 ( .in(reset_elevator2), .out(n1631) );
  inv U1370 ( .in(reset_elevator2), .out(n1632) );
  inv U1371 ( .in(reset_elevator2), .out(n1633) );
  inv U1372 ( .in(reset_elevator2), .out(n1634) );
  inv U1373 ( .in(reset_elevator2), .out(n1635) );
  inv U1374 ( .in(reset_elevator2), .out(n1636) );
  inv U1375 ( .in(reset_elevator2), .out(n1637) );
  inv U1376 ( .in(reset_elevator2), .out(n1638) );
  inv U1377 ( .in(reset_elevator2), .out(n1639) );
  inv U1378 ( .in(n1662), .out(n1640) );
  inv U1379 ( .in(n1662), .out(n1641) );
  inv U1380 ( .in(n1661), .out(n1642) );
  inv U1381 ( .in(n1661), .out(n1643) );
  inv U1382 ( .in(n1661), .out(n1644) );
  inv U1383 ( .in(n1660), .out(n1645) );
  inv U1384 ( .in(n1660), .out(n1646) );
  inv U1385 ( .in(n1660), .out(n1647) );
  inv U1386 ( .in(n1659), .out(n1648) );
  inv U1387 ( .in(n1659), .out(n1649) );
  inv U1388 ( .in(n1659), .out(n1650) );
  inv U1389 ( .in(n1658), .out(n1651) );
  inv U1390 ( .in(n1658), .out(n1652) );
  inv U1391 ( .in(n1658), .out(n1653) );
  inv U1392 ( .in(n1657), .out(n1654) );
  inv U1393 ( .in(n1657), .out(n1655) );
  inv U1394 ( .in(n1657), .out(n1656) );
  inv U1395 ( .in(reset_elevator1), .out(n1657) );
  inv U1396 ( .in(reset_elevator1), .out(n1658) );
  inv U1397 ( .in(reset_elevator1), .out(n1659) );
  inv U1398 ( .in(reset_elevator1), .out(n1660) );
  inv U1399 ( .in(reset_elevator1), .out(n1661) );
  inv U1400 ( .in(reset_elevator1), .out(n1662) );
  inv U1401 ( .in(reset_elevator1), .out(n1663) );
  inv U1402 ( .in(reset_elevator1), .out(n1664) );
  inv U1403 ( .in(reset_elevator1), .out(n1665) );
  inv U1404 ( .in(reset_elevator1), .out(n1666) );
  inv U1405 ( .in(reset_elevator1), .out(n1667) );
  inv U1406 ( .in(reset_elevator1), .out(n1668) );
  inv U1407 ( .in(reset_elevator1), .out(n1669) );
  inv U1408 ( .in(reset_elevator1), .out(n1670) );
  inv U1409 ( .in(reset_elevator1), .out(n1671) );
  inv U1410 ( .in(reset_elevator1), .out(n1672) );
  inv U1411 ( .in(reset_elevator1), .out(n1673) );
  inv U1412 ( .in(reset_elevator1), .out(n1674) );
  inv U1413 ( .in(reset_elevator1), .out(n1675) );
  inv U1414 ( .in(reset_elevator1), .out(n1676) );
  inv U1415 ( .in(reset_elevator1), .out(n1677) );
  inv U1416 ( .in(reset_elevator1), .out(n1678) );
  inv U1417 ( .in(reset_elevator1), .out(n1679) );
  inv U1418 ( .in(reset_elevator1), .out(n1680) );
  inv U1419 ( .in(reset_elevator1), .out(n1681) );
  inv U1420 ( .in(reset_elevator1), .out(n1682) );
  inv U1421 ( .in(reset_elevator1), .out(n1683) );
  inv U1422 ( .in(reset_elevator1), .out(n1684) );
  inv U1423 ( .in(final_floor_elevator2[62]), .out(n1685) );
  inv U1424 ( .in(requested_floor[62]), .out(n1686) );
  inv U1425 ( .in(n1687), .out(\ne_42/AEQB [62]) );
  inv U1426 ( .in(final_floor_elevator2[61]), .out(n1688) );
  inv U1427 ( .in(requested_floor[61]), .out(n1689) );
  inv U1428 ( .in(n1690), .out(\ne_42/AEQB [61]) );
  inv U1429 ( .in(final_floor_elevator2[60]), .out(n1691) );
  inv U1430 ( .in(requested_floor[60]), .out(n1692) );
  inv U1431 ( .in(n1693), .out(\ne_42/AEQB [60]) );
  inv U1432 ( .in(final_floor_elevator2[59]), .out(n1694) );
  inv U1433 ( .in(requested_floor[59]), .out(n1695) );
  inv U1434 ( .in(n1696), .out(\ne_42/AEQB [59]) );
  inv U1435 ( .in(final_floor_elevator2[58]), .out(n1697) );
  inv U1436 ( .in(requested_floor[58]), .out(n1698) );
  inv U1437 ( .in(n1699), .out(\ne_42/AEQB [58]) );
  inv U1438 ( .in(final_floor_elevator2[57]), .out(n1700) );
  inv U1439 ( .in(requested_floor[57]), .out(n1701) );
  inv U1440 ( .in(n1702), .out(\ne_42/AEQB [57]) );
  inv U1441 ( .in(final_floor_elevator2[56]), .out(n1703) );
  inv U1442 ( .in(requested_floor[56]), .out(n1704) );
  inv U1443 ( .in(n1705), .out(\ne_42/AEQB [56]) );
  inv U1444 ( .in(final_floor_elevator2[55]), .out(n1706) );
  inv U1445 ( .in(requested_floor[55]), .out(n1707) );
  inv U1446 ( .in(n1708), .out(\ne_42/AEQB [55]) );
  inv U1447 ( .in(final_floor_elevator2[54]), .out(n1709) );
  inv U1448 ( .in(requested_floor[54]), .out(n1710) );
  inv U1449 ( .in(n1711), .out(\ne_42/AEQB [54]) );
  inv U1450 ( .in(final_floor_elevator2[53]), .out(n1712) );
  inv U1451 ( .in(requested_floor[53]), .out(n1713) );
  inv U1452 ( .in(n1714), .out(\ne_42/AEQB [53]) );
  inv U1453 ( .in(final_floor_elevator2[52]), .out(n1715) );
  inv U1454 ( .in(requested_floor[52]), .out(n1716) );
  inv U1455 ( .in(n1717), .out(\ne_42/AEQB [52]) );
  inv U1456 ( .in(final_floor_elevator2[51]), .out(n1718) );
  inv U1457 ( .in(requested_floor[51]), .out(n1719) );
  inv U1458 ( .in(n1720), .out(\ne_42/AEQB [51]) );
  inv U1459 ( .in(final_floor_elevator2[50]), .out(n1721) );
  inv U1460 ( .in(requested_floor[50]), .out(n1722) );
  inv U1461 ( .in(n1723), .out(\ne_42/AEQB [50]) );
  inv U1462 ( .in(final_floor_elevator2[49]), .out(n1724) );
  inv U1463 ( .in(requested_floor[49]), .out(n1725) );
  inv U1464 ( .in(n1726), .out(\ne_42/AEQB [49]) );
  inv U1465 ( .in(final_floor_elevator2[48]), .out(n1727) );
  inv U1466 ( .in(requested_floor[48]), .out(n1728) );
  inv U1467 ( .in(n1729), .out(\ne_42/AEQB [48]) );
  inv U1468 ( .in(final_floor_elevator2[47]), .out(n1730) );
  inv U1469 ( .in(requested_floor[47]), .out(n1731) );
  inv U1470 ( .in(n1732), .out(\ne_42/AEQB [47]) );
  inv U1471 ( .in(final_floor_elevator2[46]), .out(n1733) );
  inv U1472 ( .in(requested_floor[46]), .out(n1734) );
  inv U1473 ( .in(n1735), .out(\ne_42/AEQB [46]) );
  inv U1474 ( .in(final_floor_elevator2[45]), .out(n1736) );
  inv U1475 ( .in(requested_floor[45]), .out(n1737) );
  inv U1476 ( .in(n1738), .out(\ne_42/AEQB [45]) );
  inv U1477 ( .in(final_floor_elevator2[44]), .out(n1739) );
  inv U1478 ( .in(requested_floor[44]), .out(n1740) );
  inv U1479 ( .in(n1741), .out(\ne_42/AEQB [44]) );
  inv U1480 ( .in(final_floor_elevator2[43]), .out(n1742) );
  inv U1481 ( .in(requested_floor[43]), .out(n1743) );
  inv U1482 ( .in(n1744), .out(\ne_42/AEQB [43]) );
  inv U1483 ( .in(final_floor_elevator2[42]), .out(n1745) );
  inv U1484 ( .in(requested_floor[42]), .out(n1746) );
  inv U1485 ( .in(n1747), .out(\ne_42/AEQB [42]) );
  inv U1486 ( .in(final_floor_elevator2[41]), .out(n1748) );
  inv U1487 ( .in(requested_floor[41]), .out(n1749) );
  inv U1488 ( .in(n1750), .out(\ne_42/AEQB [41]) );
  inv U1489 ( .in(final_floor_elevator2[40]), .out(n1751) );
  inv U1490 ( .in(requested_floor[40]), .out(n1752) );
  inv U1491 ( .in(n1753), .out(\ne_42/AEQB [40]) );
  inv U1492 ( .in(final_floor_elevator2[39]), .out(n1754) );
  inv U1493 ( .in(requested_floor[39]), .out(n1755) );
  inv U1494 ( .in(n1756), .out(\ne_42/AEQB [39]) );
  inv U1495 ( .in(final_floor_elevator2[38]), .out(n1757) );
  inv U1496 ( .in(requested_floor[38]), .out(n1758) );
  inv U1497 ( .in(n1759), .out(\ne_42/AEQB [38]) );
  inv U1498 ( .in(final_floor_elevator2[37]), .out(n1760) );
  inv U1499 ( .in(requested_floor[37]), .out(n1761) );
  inv U1500 ( .in(n1762), .out(\ne_42/AEQB [37]) );
  inv U1501 ( .in(final_floor_elevator2[36]), .out(n1763) );
  inv U1502 ( .in(requested_floor[36]), .out(n1764) );
  inv U1503 ( .in(n1765), .out(\ne_42/AEQB [36]) );
  inv U1504 ( .in(final_floor_elevator2[35]), .out(n1766) );
  inv U1505 ( .in(requested_floor[35]), .out(n1767) );
  inv U1506 ( .in(n1768), .out(\ne_42/AEQB [35]) );
  inv U1507 ( .in(final_floor_elevator2[34]), .out(n1769) );
  inv U1508 ( .in(requested_floor[34]), .out(n1770) );
  inv U1509 ( .in(n1771), .out(\ne_42/AEQB [34]) );
  inv U1510 ( .in(final_floor_elevator2[33]), .out(n1772) );
  inv U1511 ( .in(requested_floor[33]), .out(n1773) );
  inv U1512 ( .in(n1774), .out(\ne_42/AEQB [33]) );
  inv U1513 ( .in(final_floor_elevator2[32]), .out(n1775) );
  inv U1514 ( .in(requested_floor[32]), .out(n1776) );
  inv U1515 ( .in(n1777), .out(\ne_42/AEQB [32]) );
  inv U1516 ( .in(final_floor_elevator2[31]), .out(n1778) );
  inv U1517 ( .in(requested_floor[31]), .out(n1779) );
  inv U1518 ( .in(n1780), .out(\ne_42/AEQB [31]) );
  inv U1519 ( .in(final_floor_elevator2[30]), .out(n1781) );
  inv U1520 ( .in(requested_floor[30]), .out(n1782) );
  inv U1521 ( .in(n1783), .out(\ne_42/AEQB [30]) );
  inv U1522 ( .in(final_floor_elevator2[29]), .out(n1784) );
  inv U1523 ( .in(requested_floor[29]), .out(n1785) );
  inv U1524 ( .in(n1786), .out(\ne_42/AEQB [29]) );
  inv U1525 ( .in(final_floor_elevator2[28]), .out(n1787) );
  inv U1526 ( .in(requested_floor[28]), .out(n1788) );
  inv U1527 ( .in(n1789), .out(\ne_42/AEQB [28]) );
  inv U1528 ( .in(final_floor_elevator2[27]), .out(n1790) );
  inv U1529 ( .in(requested_floor[27]), .out(n1791) );
  inv U1530 ( .in(n1792), .out(\ne_42/AEQB [27]) );
  inv U1531 ( .in(final_floor_elevator2[26]), .out(n1793) );
  inv U1532 ( .in(requested_floor[26]), .out(n1794) );
  inv U1533 ( .in(n1795), .out(\ne_42/AEQB [26]) );
  inv U1534 ( .in(final_floor_elevator2[25]), .out(n1796) );
  inv U1535 ( .in(requested_floor[25]), .out(n1797) );
  inv U1536 ( .in(n1798), .out(\ne_42/AEQB [25]) );
  inv U1537 ( .in(final_floor_elevator2[24]), .out(n1799) );
  inv U1538 ( .in(requested_floor[24]), .out(n1800) );
  inv U1539 ( .in(n1801), .out(\ne_42/AEQB [24]) );
  inv U1540 ( .in(final_floor_elevator2[23]), .out(n1802) );
  inv U1541 ( .in(requested_floor[23]), .out(n1803) );
  inv U1542 ( .in(n1804), .out(\ne_42/AEQB [23]) );
  inv U1543 ( .in(final_floor_elevator2[22]), .out(n1805) );
  inv U1544 ( .in(requested_floor[22]), .out(n1806) );
  inv U1545 ( .in(n1807), .out(\ne_42/AEQB [22]) );
  inv U1546 ( .in(final_floor_elevator2[21]), .out(n1808) );
  inv U1547 ( .in(requested_floor[21]), .out(n1809) );
  inv U1548 ( .in(n1810), .out(\ne_42/AEQB [21]) );
  inv U1549 ( .in(final_floor_elevator2[20]), .out(n1811) );
  inv U1550 ( .in(requested_floor[20]), .out(n1812) );
  inv U1551 ( .in(n1813), .out(\ne_42/AEQB [20]) );
  inv U1552 ( .in(final_floor_elevator2[19]), .out(n1814) );
  inv U1553 ( .in(requested_floor[19]), .out(n1815) );
  inv U1554 ( .in(n1816), .out(\ne_42/AEQB [19]) );
  inv U1555 ( .in(final_floor_elevator2[18]), .out(n1817) );
  inv U1556 ( .in(requested_floor[18]), .out(n1818) );
  inv U1557 ( .in(n1819), .out(\ne_42/AEQB [18]) );
  inv U1558 ( .in(final_floor_elevator2[17]), .out(n1820) );
  inv U1559 ( .in(requested_floor[17]), .out(n1821) );
  inv U1560 ( .in(n1822), .out(\ne_42/AEQB [17]) );
  inv U1561 ( .in(final_floor_elevator2[16]), .out(n1823) );
  inv U1562 ( .in(requested_floor[16]), .out(n1824) );
  inv U1563 ( .in(n1825), .out(\ne_42/AEQB [16]) );
  inv U1564 ( .in(final_floor_elevator2[15]), .out(n1826) );
  inv U1565 ( .in(requested_floor[15]), .out(n1827) );
  inv U1566 ( .in(n1828), .out(\ne_42/AEQB [15]) );
  inv U1567 ( .in(final_floor_elevator2[14]), .out(n1829) );
  inv U1568 ( .in(requested_floor[14]), .out(n1830) );
  inv U1569 ( .in(n1831), .out(\ne_42/AEQB [14]) );
  inv U1570 ( .in(final_floor_elevator2[13]), .out(n1832) );
  inv U1571 ( .in(requested_floor[13]), .out(n1833) );
  inv U1572 ( .in(n1834), .out(\ne_42/AEQB [13]) );
  inv U1573 ( .in(final_floor_elevator2[12]), .out(n1835) );
  inv U1574 ( .in(requested_floor[12]), .out(n1836) );
  inv U1575 ( .in(n1837), .out(\ne_42/AEQB [12]) );
  inv U1576 ( .in(final_floor_elevator2[11]), .out(n1838) );
  inv U1577 ( .in(requested_floor[11]), .out(n1839) );
  inv U1578 ( .in(n1840), .out(\ne_42/AEQB [11]) );
  inv U1579 ( .in(final_floor_elevator2[10]), .out(n1841) );
  inv U1580 ( .in(requested_floor[10]), .out(n1842) );
  inv U1581 ( .in(n1843), .out(\ne_42/AEQB [10]) );
  inv U1582 ( .in(final_floor_elevator2[9]), .out(n1844) );
  inv U1583 ( .in(requested_floor[9]), .out(n1845) );
  inv U1584 ( .in(n1846), .out(\ne_42/AEQB [9]) );
  inv U1585 ( .in(final_floor_elevator2[8]), .out(n1847) );
  inv U1586 ( .in(requested_floor[8]), .out(n1848) );
  inv U1587 ( .in(n1849), .out(\ne_42/AEQB [8]) );
  inv U1588 ( .in(final_floor_elevator2[7]), .out(n1850) );
  inv U1589 ( .in(requested_floor[7]), .out(n1851) );
  inv U1590 ( .in(n1852), .out(\ne_42/AEQB [7]) );
  inv U1591 ( .in(final_floor_elevator2[6]), .out(n1853) );
  inv U1592 ( .in(requested_floor[6]), .out(n1854) );
  inv U1593 ( .in(n1855), .out(\ne_42/AEQB [6]) );
  inv U1594 ( .in(final_floor_elevator2[5]), .out(n1856) );
  inv U1595 ( .in(requested_floor[5]), .out(n1857) );
  inv U1596 ( .in(n1858), .out(\ne_42/AEQB [5]) );
  inv U1597 ( .in(final_floor_elevator2[4]), .out(n1859) );
  inv U1598 ( .in(requested_floor[4]), .out(n1860) );
  inv U1599 ( .in(n1861), .out(\ne_42/AEQB [4]) );
  inv U1600 ( .in(final_floor_elevator2[3]), .out(n1862) );
  inv U1601 ( .in(requested_floor[3]), .out(n1863) );
  inv U1602 ( .in(n1864), .out(\ne_42/AEQB [3]) );
  inv U1603 ( .in(final_floor_elevator2[2]), .out(n1865) );
  inv U1604 ( .in(requested_floor[2]), .out(n1866) );
  inv U1605 ( .in(n1867), .out(\ne_42/AEQB [2]) );
  inv U1606 ( .in(final_floor_elevator2[1]), .out(n1868) );
  inv U1607 ( .in(requested_floor[1]), .out(n1869) );
  inv U1608 ( .in(n1870), .out(\ne_42/AEQB [1]) );
  inv U1609 ( .in(\ne_42/SA ), .out(n1871) );
  inv U1610 ( .in(\ne_47/SB ), .out(n1872) );
  inv U1611 ( .in(n1873), .out(\ne_42/AEQB [63]) );
  inv U1612 ( .in(n1874), .out(\ne_42/LTV [1]) );
  inv U1613 ( .in(final_floor_elevator2[0]), .out(n1875) );
  inv U1614 ( .in(n1876), .out(\ne_42/GTV [1]) );
  inv U1615 ( .in(requested_floor[0]), .out(n1877) );
  inv U1616 ( .in(current_floor_output_elevator1[62]), .out(n1878) );
  inv U1617 ( .in(destination_floor_elevator1[62]), .out(n1879) );
  inv U1618 ( .in(n1880), .out(\eq_42_3/AEQB [62]) );
  inv U1619 ( .in(current_floor_output_elevator1[61]), .out(n1881) );
  inv U1620 ( .in(destination_floor_elevator1[61]), .out(n1882) );
  inv U1621 ( .in(n1883), .out(\eq_42_3/AEQB [61]) );
  inv U1622 ( .in(current_floor_output_elevator1[60]), .out(n1884) );
  inv U1623 ( .in(destination_floor_elevator1[60]), .out(n1885) );
  inv U1624 ( .in(n1886), .out(\eq_42_3/AEQB [60]) );
  inv U1625 ( .in(current_floor_output_elevator1[59]), .out(n1887) );
  inv U1626 ( .in(destination_floor_elevator1[59]), .out(n1888) );
  inv U1627 ( .in(n1889), .out(\eq_42_3/AEQB [59]) );
  inv U1628 ( .in(current_floor_output_elevator1[58]), .out(n1890) );
  inv U1629 ( .in(destination_floor_elevator1[58]), .out(n1891) );
  inv U1630 ( .in(n1892), .out(\eq_42_3/AEQB [58]) );
  inv U1631 ( .in(current_floor_output_elevator1[57]), .out(n1893) );
  inv U1632 ( .in(destination_floor_elevator1[57]), .out(n1894) );
  inv U1633 ( .in(n1895), .out(\eq_42_3/AEQB [57]) );
  inv U1634 ( .in(current_floor_output_elevator1[56]), .out(n1896) );
  inv U1635 ( .in(destination_floor_elevator1[56]), .out(n1897) );
  inv U1636 ( .in(n1898), .out(\eq_42_3/AEQB [56]) );
  inv U1637 ( .in(current_floor_output_elevator1[55]), .out(n1899) );
  inv U1638 ( .in(destination_floor_elevator1[55]), .out(n1900) );
  inv U1639 ( .in(n1901), .out(\eq_42_3/AEQB [55]) );
  inv U1640 ( .in(current_floor_output_elevator1[54]), .out(n1902) );
  inv U1641 ( .in(destination_floor_elevator1[54]), .out(n1903) );
  inv U1642 ( .in(n1904), .out(\eq_42_3/AEQB [54]) );
  inv U1643 ( .in(current_floor_output_elevator1[53]), .out(n1905) );
  inv U1644 ( .in(destination_floor_elevator1[53]), .out(n1906) );
  inv U1645 ( .in(n1907), .out(\eq_42_3/AEQB [53]) );
  inv U1646 ( .in(current_floor_output_elevator1[52]), .out(n1908) );
  inv U1647 ( .in(destination_floor_elevator1[52]), .out(n1909) );
  inv U1648 ( .in(n1910), .out(\eq_42_3/AEQB [52]) );
  inv U1649 ( .in(current_floor_output_elevator1[51]), .out(n1911) );
  inv U1650 ( .in(destination_floor_elevator1[51]), .out(n1912) );
  inv U1651 ( .in(n1913), .out(\eq_42_3/AEQB [51]) );
  inv U1652 ( .in(current_floor_output_elevator1[50]), .out(n1914) );
  inv U1653 ( .in(destination_floor_elevator1[50]), .out(n1915) );
  inv U1654 ( .in(n1916), .out(\eq_42_3/AEQB [50]) );
  inv U1655 ( .in(current_floor_output_elevator1[49]), .out(n1917) );
  inv U1656 ( .in(destination_floor_elevator1[49]), .out(n1918) );
  inv U1657 ( .in(n1919), .out(\eq_42_3/AEQB [49]) );
  inv U1658 ( .in(current_floor_output_elevator1[48]), .out(n1920) );
  inv U1659 ( .in(destination_floor_elevator1[48]), .out(n1921) );
  inv U1660 ( .in(n1922), .out(\eq_42_3/AEQB [48]) );
  inv U1661 ( .in(current_floor_output_elevator1[47]), .out(n1923) );
  inv U1662 ( .in(destination_floor_elevator1[47]), .out(n1924) );
  inv U1663 ( .in(n1925), .out(\eq_42_3/AEQB [47]) );
  inv U1664 ( .in(current_floor_output_elevator1[46]), .out(n1926) );
  inv U1665 ( .in(destination_floor_elevator1[46]), .out(n1927) );
  inv U1666 ( .in(n1928), .out(\eq_42_3/AEQB [46]) );
  inv U1667 ( .in(current_floor_output_elevator1[45]), .out(n1929) );
  inv U1668 ( .in(destination_floor_elevator1[45]), .out(n1930) );
  inv U1669 ( .in(n1931), .out(\eq_42_3/AEQB [45]) );
  inv U1670 ( .in(current_floor_output_elevator1[44]), .out(n1932) );
  inv U1671 ( .in(destination_floor_elevator1[44]), .out(n1933) );
  inv U1672 ( .in(n1934), .out(\eq_42_3/AEQB [44]) );
  inv U1673 ( .in(current_floor_output_elevator1[43]), .out(n1935) );
  inv U1674 ( .in(destination_floor_elevator1[43]), .out(n1936) );
  inv U1675 ( .in(n1937), .out(\eq_42_3/AEQB [43]) );
  inv U1676 ( .in(current_floor_output_elevator1[42]), .out(n1938) );
  inv U1677 ( .in(destination_floor_elevator1[42]), .out(n1939) );
  inv U1678 ( .in(n1940), .out(\eq_42_3/AEQB [42]) );
  inv U1679 ( .in(current_floor_output_elevator1[41]), .out(n1941) );
  inv U1680 ( .in(destination_floor_elevator1[41]), .out(n1942) );
  inv U1681 ( .in(n1943), .out(\eq_42_3/AEQB [41]) );
  inv U1682 ( .in(current_floor_output_elevator1[40]), .out(n1944) );
  inv U1683 ( .in(destination_floor_elevator1[40]), .out(n1945) );
  inv U1684 ( .in(n1946), .out(\eq_42_3/AEQB [40]) );
  inv U1685 ( .in(current_floor_output_elevator1[39]), .out(n1947) );
  inv U1686 ( .in(destination_floor_elevator1[39]), .out(n1948) );
  inv U1687 ( .in(n1949), .out(\eq_42_3/AEQB [39]) );
  inv U1688 ( .in(current_floor_output_elevator1[38]), .out(n1950) );
  inv U1689 ( .in(destination_floor_elevator1[38]), .out(n1951) );
  inv U1690 ( .in(n1952), .out(\eq_42_3/AEQB [38]) );
  inv U1691 ( .in(current_floor_output_elevator1[37]), .out(n1953) );
  inv U1692 ( .in(destination_floor_elevator1[37]), .out(n1954) );
  inv U1693 ( .in(n1955), .out(\eq_42_3/AEQB [37]) );
  inv U1694 ( .in(current_floor_output_elevator1[36]), .out(n1956) );
  inv U1695 ( .in(destination_floor_elevator1[36]), .out(n1957) );
  inv U1696 ( .in(n1958), .out(\eq_42_3/AEQB [36]) );
  inv U1697 ( .in(current_floor_output_elevator1[35]), .out(n1959) );
  inv U1698 ( .in(destination_floor_elevator1[35]), .out(n1960) );
  inv U1699 ( .in(n1961), .out(\eq_42_3/AEQB [35]) );
  inv U1700 ( .in(current_floor_output_elevator1[34]), .out(n1962) );
  inv U1701 ( .in(destination_floor_elevator1[34]), .out(n1963) );
  inv U1702 ( .in(n1964), .out(\eq_42_3/AEQB [34]) );
  inv U1703 ( .in(current_floor_output_elevator1[33]), .out(n1965) );
  inv U1704 ( .in(destination_floor_elevator1[33]), .out(n1966) );
  inv U1705 ( .in(n1967), .out(\eq_42_3/AEQB [33]) );
  inv U1706 ( .in(current_floor_output_elevator1[32]), .out(n1968) );
  inv U1707 ( .in(destination_floor_elevator1[32]), .out(n1969) );
  inv U1708 ( .in(n1970), .out(\eq_42_3/AEQB [32]) );
  inv U1709 ( .in(current_floor_output_elevator1[31]), .out(n1971) );
  inv U1710 ( .in(destination_floor_elevator1[31]), .out(n1972) );
  inv U1711 ( .in(n1973), .out(\eq_42_3/AEQB [31]) );
  inv U1712 ( .in(current_floor_output_elevator1[30]), .out(n1974) );
  inv U1713 ( .in(destination_floor_elevator1[30]), .out(n1975) );
  inv U1714 ( .in(n1976), .out(\eq_42_3/AEQB [30]) );
  inv U1715 ( .in(current_floor_output_elevator1[29]), .out(n1977) );
  inv U1716 ( .in(destination_floor_elevator1[29]), .out(n1978) );
  inv U1717 ( .in(n1979), .out(\eq_42_3/AEQB [29]) );
  inv U1718 ( .in(current_floor_output_elevator1[28]), .out(n1980) );
  inv U1719 ( .in(destination_floor_elevator1[28]), .out(n1981) );
  inv U1720 ( .in(n1982), .out(\eq_42_3/AEQB [28]) );
  inv U1721 ( .in(current_floor_output_elevator1[27]), .out(n1983) );
  inv U1722 ( .in(destination_floor_elevator1[27]), .out(n1984) );
  inv U1723 ( .in(n1985), .out(\eq_42_3/AEQB [27]) );
  inv U1724 ( .in(current_floor_output_elevator1[26]), .out(n1986) );
  inv U1725 ( .in(destination_floor_elevator1[26]), .out(n1987) );
  inv U1726 ( .in(n1988), .out(\eq_42_3/AEQB [26]) );
  inv U1727 ( .in(current_floor_output_elevator1[25]), .out(n1989) );
  inv U1728 ( .in(destination_floor_elevator1[25]), .out(n1990) );
  inv U1729 ( .in(n1991), .out(\eq_42_3/AEQB [25]) );
  inv U1730 ( .in(current_floor_output_elevator1[24]), .out(n1992) );
  inv U1731 ( .in(destination_floor_elevator1[24]), .out(n1993) );
  inv U1732 ( .in(n1994), .out(\eq_42_3/AEQB [24]) );
  inv U1733 ( .in(current_floor_output_elevator1[23]), .out(n1995) );
  inv U1734 ( .in(destination_floor_elevator1[23]), .out(n1996) );
  inv U1735 ( .in(n1997), .out(\eq_42_3/AEQB [23]) );
  inv U1736 ( .in(current_floor_output_elevator1[22]), .out(n1998) );
  inv U1737 ( .in(destination_floor_elevator1[22]), .out(n1999) );
  inv U1738 ( .in(n2000), .out(\eq_42_3/AEQB [22]) );
  inv U1739 ( .in(current_floor_output_elevator1[21]), .out(n2001) );
  inv U1740 ( .in(destination_floor_elevator1[21]), .out(n2002) );
  inv U1741 ( .in(n2003), .out(\eq_42_3/AEQB [21]) );
  inv U1742 ( .in(current_floor_output_elevator1[20]), .out(n2004) );
  inv U1743 ( .in(destination_floor_elevator1[20]), .out(n2005) );
  inv U1744 ( .in(n2006), .out(\eq_42_3/AEQB [20]) );
  inv U1745 ( .in(current_floor_output_elevator1[19]), .out(n2007) );
  inv U1746 ( .in(destination_floor_elevator1[19]), .out(n2008) );
  inv U1747 ( .in(n2009), .out(\eq_42_3/AEQB [19]) );
  inv U1748 ( .in(current_floor_output_elevator1[18]), .out(n2010) );
  inv U1749 ( .in(destination_floor_elevator1[18]), .out(n2011) );
  inv U1750 ( .in(n2012), .out(\eq_42_3/AEQB [18]) );
  inv U1751 ( .in(current_floor_output_elevator1[17]), .out(n2013) );
  inv U1752 ( .in(destination_floor_elevator1[17]), .out(n2014) );
  inv U1753 ( .in(n2015), .out(\eq_42_3/AEQB [17]) );
  inv U1754 ( .in(current_floor_output_elevator1[16]), .out(n2016) );
  inv U1755 ( .in(destination_floor_elevator1[16]), .out(n2017) );
  inv U1756 ( .in(n2018), .out(\eq_42_3/AEQB [16]) );
  inv U1757 ( .in(current_floor_output_elevator1[15]), .out(n2019) );
  inv U1758 ( .in(destination_floor_elevator1[15]), .out(n2020) );
  inv U1759 ( .in(n2021), .out(\eq_42_3/AEQB [15]) );
  inv U1760 ( .in(current_floor_output_elevator1[14]), .out(n2022) );
  inv U1761 ( .in(destination_floor_elevator1[14]), .out(n2023) );
  inv U1762 ( .in(n2024), .out(\eq_42_3/AEQB [14]) );
  inv U1763 ( .in(current_floor_output_elevator1[13]), .out(n2025) );
  inv U1764 ( .in(destination_floor_elevator1[13]), .out(n2026) );
  inv U1765 ( .in(n2027), .out(\eq_42_3/AEQB [13]) );
  inv U1766 ( .in(current_floor_output_elevator1[12]), .out(n2028) );
  inv U1767 ( .in(destination_floor_elevator1[12]), .out(n2029) );
  inv U1768 ( .in(n2030), .out(\eq_42_3/AEQB [12]) );
  inv U1769 ( .in(current_floor_output_elevator1[11]), .out(n2031) );
  inv U1770 ( .in(destination_floor_elevator1[11]), .out(n2032) );
  inv U1771 ( .in(n2033), .out(\eq_42_3/AEQB [11]) );
  inv U1772 ( .in(current_floor_output_elevator1[10]), .out(n2034) );
  inv U1773 ( .in(destination_floor_elevator1[10]), .out(n2035) );
  inv U1774 ( .in(n2036), .out(\eq_42_3/AEQB [10]) );
  inv U1775 ( .in(current_floor_output_elevator1[9]), .out(n2037) );
  inv U1776 ( .in(destination_floor_elevator1[9]), .out(n2038) );
  inv U1777 ( .in(n2039), .out(\eq_42_3/AEQB [9]) );
  inv U1778 ( .in(current_floor_output_elevator1[8]), .out(n2040) );
  inv U1779 ( .in(destination_floor_elevator1[8]), .out(n2041) );
  inv U1780 ( .in(n2042), .out(\eq_42_3/AEQB [8]) );
  inv U1781 ( .in(current_floor_output_elevator1[7]), .out(n2043) );
  inv U1782 ( .in(destination_floor_elevator1[7]), .out(n2044) );
  inv U1783 ( .in(n2045), .out(\eq_42_3/AEQB [7]) );
  inv U1784 ( .in(current_floor_output_elevator1[6]), .out(n2046) );
  inv U1785 ( .in(destination_floor_elevator1[6]), .out(n2047) );
  inv U1786 ( .in(n2048), .out(\eq_42_3/AEQB [6]) );
  inv U1787 ( .in(current_floor_output_elevator1[5]), .out(n2049) );
  inv U1788 ( .in(destination_floor_elevator1[5]), .out(n2050) );
  inv U1789 ( .in(n2051), .out(\eq_42_3/AEQB [5]) );
  inv U1790 ( .in(current_floor_output_elevator1[4]), .out(n2052) );
  inv U1791 ( .in(destination_floor_elevator1[4]), .out(n2053) );
  inv U1792 ( .in(n2054), .out(\eq_42_3/AEQB [4]) );
  inv U1793 ( .in(current_floor_output_elevator1[3]), .out(n2055) );
  inv U1794 ( .in(destination_floor_elevator1[3]), .out(n2056) );
  inv U1795 ( .in(n2057), .out(\eq_42_3/AEQB [3]) );
  inv U1796 ( .in(current_floor_output_elevator1[2]), .out(n2058) );
  inv U1797 ( .in(destination_floor_elevator1[2]), .out(n2059) );
  inv U1798 ( .in(n2060), .out(\eq_42_3/AEQB [2]) );
  inv U1799 ( .in(current_floor_output_elevator1[1]), .out(n2061) );
  inv U1800 ( .in(destination_floor_elevator1[1]), .out(n2062) );
  inv U1801 ( .in(n2063), .out(\eq_42_3/AEQB [1]) );
  inv U1802 ( .in(\eq_42_3/SA ), .out(n2064) );
  inv U1803 ( .in(\eq_42_3/SB ), .out(n2065) );
  inv U1804 ( .in(n2066), .out(\eq_42_3/AEQB [63]) );
  inv U1805 ( .in(n2067), .out(\eq_42_3/LTV [1]) );
  inv U1806 ( .in(current_floor_output_elevator1[0]), .out(n2068) );
  inv U1807 ( .in(n2069), .out(\eq_42_3/GTV [1]) );
  inv U1808 ( .in(destination_floor_elevator1[0]), .out(n2070) );
  inv U1809 ( .in(final_floor_elevator1[62]), .out(n2071) );
  inv U1810 ( .in(requested_floor[62]), .out(n2072) );
  inv U1811 ( .in(n2073), .out(\ne_47/AEQB [62]) );
  inv U1812 ( .in(final_floor_elevator1[61]), .out(n2074) );
  inv U1813 ( .in(requested_floor[61]), .out(n2075) );
  inv U1814 ( .in(n2076), .out(\ne_47/AEQB [61]) );
  inv U1815 ( .in(final_floor_elevator1[60]), .out(n2077) );
  inv U1816 ( .in(requested_floor[60]), .out(n2078) );
  inv U1817 ( .in(n2079), .out(\ne_47/AEQB [60]) );
  inv U1818 ( .in(final_floor_elevator1[59]), .out(n2080) );
  inv U1819 ( .in(requested_floor[59]), .out(n2081) );
  inv U1820 ( .in(n2082), .out(\ne_47/AEQB [59]) );
  inv U1821 ( .in(final_floor_elevator1[58]), .out(n2083) );
  inv U1822 ( .in(requested_floor[58]), .out(n2084) );
  inv U1823 ( .in(n2085), .out(\ne_47/AEQB [58]) );
  inv U1824 ( .in(final_floor_elevator1[57]), .out(n2086) );
  inv U1825 ( .in(requested_floor[57]), .out(n2087) );
  inv U1826 ( .in(n2088), .out(\ne_47/AEQB [57]) );
  inv U1827 ( .in(final_floor_elevator1[56]), .out(n2089) );
  inv U1828 ( .in(requested_floor[56]), .out(n2090) );
  inv U1829 ( .in(n2091), .out(\ne_47/AEQB [56]) );
  inv U1830 ( .in(final_floor_elevator1[55]), .out(n2092) );
  inv U1831 ( .in(requested_floor[55]), .out(n2093) );
  inv U1832 ( .in(n2094), .out(\ne_47/AEQB [55]) );
  inv U1833 ( .in(final_floor_elevator1[54]), .out(n2095) );
  inv U1834 ( .in(requested_floor[54]), .out(n2096) );
  inv U1835 ( .in(n2097), .out(\ne_47/AEQB [54]) );
  inv U1836 ( .in(final_floor_elevator1[53]), .out(n2098) );
  inv U1837 ( .in(requested_floor[53]), .out(n2099) );
  inv U1838 ( .in(n2100), .out(\ne_47/AEQB [53]) );
  inv U1839 ( .in(final_floor_elevator1[52]), .out(n2101) );
  inv U1840 ( .in(requested_floor[52]), .out(n2102) );
  inv U1841 ( .in(n2103), .out(\ne_47/AEQB [52]) );
  inv U1842 ( .in(final_floor_elevator1[51]), .out(n2104) );
  inv U1843 ( .in(requested_floor[51]), .out(n2105) );
  inv U1844 ( .in(n2106), .out(\ne_47/AEQB [51]) );
  inv U1845 ( .in(final_floor_elevator1[50]), .out(n2107) );
  inv U1846 ( .in(requested_floor[50]), .out(n2108) );
  inv U1847 ( .in(n2109), .out(\ne_47/AEQB [50]) );
  inv U1848 ( .in(final_floor_elevator1[49]), .out(n2110) );
  inv U1849 ( .in(requested_floor[49]), .out(n2111) );
  inv U1850 ( .in(n2112), .out(\ne_47/AEQB [49]) );
  inv U1851 ( .in(final_floor_elevator1[48]), .out(n2113) );
  inv U1852 ( .in(requested_floor[48]), .out(n2114) );
  inv U1853 ( .in(n2115), .out(\ne_47/AEQB [48]) );
  inv U1854 ( .in(final_floor_elevator1[47]), .out(n2116) );
  inv U1855 ( .in(requested_floor[47]), .out(n2117) );
  inv U1856 ( .in(n2118), .out(\ne_47/AEQB [47]) );
  inv U1857 ( .in(final_floor_elevator1[46]), .out(n2119) );
  inv U1858 ( .in(requested_floor[46]), .out(n2120) );
  inv U1859 ( .in(n2121), .out(\ne_47/AEQB [46]) );
  inv U1860 ( .in(final_floor_elevator1[45]), .out(n2122) );
  inv U1861 ( .in(requested_floor[45]), .out(n2123) );
  inv U1862 ( .in(n2124), .out(\ne_47/AEQB [45]) );
  inv U1863 ( .in(final_floor_elevator1[44]), .out(n2125) );
  inv U1864 ( .in(requested_floor[44]), .out(n2126) );
  inv U1865 ( .in(n2127), .out(\ne_47/AEQB [44]) );
  inv U1866 ( .in(final_floor_elevator1[43]), .out(n2128) );
  inv U1867 ( .in(requested_floor[43]), .out(n2129) );
  inv U1868 ( .in(n2130), .out(\ne_47/AEQB [43]) );
  inv U1869 ( .in(final_floor_elevator1[42]), .out(n2131) );
  inv U1870 ( .in(requested_floor[42]), .out(n2132) );
  inv U1871 ( .in(n2133), .out(\ne_47/AEQB [42]) );
  inv U1872 ( .in(final_floor_elevator1[41]), .out(n2134) );
  inv U1873 ( .in(requested_floor[41]), .out(n2135) );
  inv U1874 ( .in(n2136), .out(\ne_47/AEQB [41]) );
  inv U1875 ( .in(final_floor_elevator1[40]), .out(n2137) );
  inv U1876 ( .in(requested_floor[40]), .out(n2138) );
  inv U1877 ( .in(n2139), .out(\ne_47/AEQB [40]) );
  inv U1878 ( .in(final_floor_elevator1[39]), .out(n2140) );
  inv U1879 ( .in(requested_floor[39]), .out(n2141) );
  inv U1880 ( .in(n2142), .out(\ne_47/AEQB [39]) );
  inv U1881 ( .in(final_floor_elevator1[38]), .out(n2143) );
  inv U1882 ( .in(requested_floor[38]), .out(n2144) );
  inv U1883 ( .in(n2145), .out(\ne_47/AEQB [38]) );
  inv U1884 ( .in(final_floor_elevator1[37]), .out(n2146) );
  inv U1885 ( .in(requested_floor[37]), .out(n2147) );
  inv U1886 ( .in(n2148), .out(\ne_47/AEQB [37]) );
  inv U1887 ( .in(final_floor_elevator1[36]), .out(n2149) );
  inv U1888 ( .in(requested_floor[36]), .out(n2150) );
  inv U1889 ( .in(n2151), .out(\ne_47/AEQB [36]) );
  inv U1890 ( .in(final_floor_elevator1[35]), .out(n2152) );
  inv U1891 ( .in(requested_floor[35]), .out(n2153) );
  inv U1892 ( .in(n2154), .out(\ne_47/AEQB [35]) );
  inv U1893 ( .in(final_floor_elevator1[34]), .out(n2155) );
  inv U1894 ( .in(requested_floor[34]), .out(n2156) );
  inv U1895 ( .in(n2157), .out(\ne_47/AEQB [34]) );
  inv U1896 ( .in(final_floor_elevator1[33]), .out(n2158) );
  inv U1897 ( .in(requested_floor[33]), .out(n2159) );
  inv U1898 ( .in(n2160), .out(\ne_47/AEQB [33]) );
  inv U1899 ( .in(final_floor_elevator1[32]), .out(n2161) );
  inv U1900 ( .in(requested_floor[32]), .out(n2162) );
  inv U1901 ( .in(n2163), .out(\ne_47/AEQB [32]) );
  inv U1902 ( .in(final_floor_elevator1[31]), .out(n2164) );
  inv U1903 ( .in(requested_floor[31]), .out(n2165) );
  inv U1904 ( .in(n2166), .out(\ne_47/AEQB [31]) );
  inv U1905 ( .in(final_floor_elevator1[30]), .out(n2167) );
  inv U1906 ( .in(requested_floor[30]), .out(n2168) );
  inv U1907 ( .in(n2169), .out(\ne_47/AEQB [30]) );
  inv U1908 ( .in(final_floor_elevator1[29]), .out(n2170) );
  inv U1909 ( .in(requested_floor[29]), .out(n2171) );
  inv U1910 ( .in(n2172), .out(\ne_47/AEQB [29]) );
  inv U1911 ( .in(final_floor_elevator1[28]), .out(n2173) );
  inv U1912 ( .in(requested_floor[28]), .out(n2174) );
  inv U1913 ( .in(n2175), .out(\ne_47/AEQB [28]) );
  inv U1914 ( .in(final_floor_elevator1[27]), .out(n2176) );
  inv U1915 ( .in(requested_floor[27]), .out(n2177) );
  inv U1916 ( .in(n2178), .out(\ne_47/AEQB [27]) );
  inv U1917 ( .in(final_floor_elevator1[26]), .out(n2179) );
  inv U1918 ( .in(requested_floor[26]), .out(n2180) );
  inv U1919 ( .in(n2181), .out(\ne_47/AEQB [26]) );
  inv U1920 ( .in(final_floor_elevator1[25]), .out(n2182) );
  inv U1921 ( .in(requested_floor[25]), .out(n2183) );
  inv U1922 ( .in(n2184), .out(\ne_47/AEQB [25]) );
  inv U1923 ( .in(final_floor_elevator1[24]), .out(n2185) );
  inv U1924 ( .in(requested_floor[24]), .out(n2186) );
  inv U1925 ( .in(n2187), .out(\ne_47/AEQB [24]) );
  inv U1926 ( .in(final_floor_elevator1[23]), .out(n2188) );
  inv U1927 ( .in(requested_floor[23]), .out(n2189) );
  inv U1928 ( .in(n2190), .out(\ne_47/AEQB [23]) );
  inv U1929 ( .in(final_floor_elevator1[22]), .out(n2191) );
  inv U1930 ( .in(requested_floor[22]), .out(n2192) );
  inv U1931 ( .in(n2193), .out(\ne_47/AEQB [22]) );
  inv U1932 ( .in(final_floor_elevator1[21]), .out(n2194) );
  inv U1933 ( .in(requested_floor[21]), .out(n2195) );
  inv U1934 ( .in(n2196), .out(\ne_47/AEQB [21]) );
  inv U1935 ( .in(final_floor_elevator1[20]), .out(n2197) );
  inv U1936 ( .in(requested_floor[20]), .out(n2198) );
  inv U1937 ( .in(n2199), .out(\ne_47/AEQB [20]) );
  inv U1938 ( .in(final_floor_elevator1[19]), .out(n2200) );
  inv U1939 ( .in(requested_floor[19]), .out(n2201) );
  inv U1940 ( .in(n2202), .out(\ne_47/AEQB [19]) );
  inv U1941 ( .in(final_floor_elevator1[18]), .out(n2203) );
  inv U1942 ( .in(requested_floor[18]), .out(n2204) );
  inv U1943 ( .in(n2205), .out(\ne_47/AEQB [18]) );
  inv U1944 ( .in(final_floor_elevator1[17]), .out(n2206) );
  inv U1945 ( .in(requested_floor[17]), .out(n2207) );
  inv U1946 ( .in(n2208), .out(\ne_47/AEQB [17]) );
  inv U1947 ( .in(final_floor_elevator1[16]), .out(n2209) );
  inv U1948 ( .in(requested_floor[16]), .out(n2210) );
  inv U1949 ( .in(n2211), .out(\ne_47/AEQB [16]) );
  inv U1950 ( .in(final_floor_elevator1[15]), .out(n2212) );
  inv U1951 ( .in(requested_floor[15]), .out(n2213) );
  inv U1952 ( .in(n2214), .out(\ne_47/AEQB [15]) );
  inv U1953 ( .in(final_floor_elevator1[14]), .out(n2215) );
  inv U1954 ( .in(requested_floor[14]), .out(n2216) );
  inv U1955 ( .in(n2217), .out(\ne_47/AEQB [14]) );
  inv U1956 ( .in(final_floor_elevator1[13]), .out(n2218) );
  inv U1957 ( .in(requested_floor[13]), .out(n2219) );
  inv U1958 ( .in(n2220), .out(\ne_47/AEQB [13]) );
  inv U1959 ( .in(final_floor_elevator1[12]), .out(n2221) );
  inv U1960 ( .in(requested_floor[12]), .out(n2222) );
  inv U1961 ( .in(n2223), .out(\ne_47/AEQB [12]) );
  inv U1962 ( .in(final_floor_elevator1[11]), .out(n2224) );
  inv U1963 ( .in(requested_floor[11]), .out(n2225) );
  inv U1964 ( .in(n2226), .out(\ne_47/AEQB [11]) );
  inv U1965 ( .in(final_floor_elevator1[10]), .out(n2227) );
  inv U1966 ( .in(requested_floor[10]), .out(n2228) );
  inv U1967 ( .in(n2229), .out(\ne_47/AEQB [10]) );
  inv U1968 ( .in(final_floor_elevator1[9]), .out(n2230) );
  inv U1969 ( .in(requested_floor[9]), .out(n2231) );
  inv U1970 ( .in(n2232), .out(\ne_47/AEQB [9]) );
  inv U1971 ( .in(final_floor_elevator1[8]), .out(n2233) );
  inv U1972 ( .in(requested_floor[8]), .out(n2234) );
  inv U1973 ( .in(n2235), .out(\ne_47/AEQB [8]) );
  inv U1974 ( .in(final_floor_elevator1[7]), .out(n2236) );
  inv U1975 ( .in(requested_floor[7]), .out(n2237) );
  inv U1976 ( .in(n2238), .out(\ne_47/AEQB [7]) );
  inv U1977 ( .in(final_floor_elevator1[6]), .out(n2239) );
  inv U1978 ( .in(requested_floor[6]), .out(n2240) );
  inv U1979 ( .in(n2241), .out(\ne_47/AEQB [6]) );
  inv U1980 ( .in(final_floor_elevator1[5]), .out(n2242) );
  inv U1981 ( .in(requested_floor[5]), .out(n2243) );
  inv U1982 ( .in(n2244), .out(\ne_47/AEQB [5]) );
  inv U1983 ( .in(final_floor_elevator1[4]), .out(n2245) );
  inv U1984 ( .in(requested_floor[4]), .out(n2246) );
  inv U1985 ( .in(n2247), .out(\ne_47/AEQB [4]) );
  inv U1986 ( .in(final_floor_elevator1[3]), .out(n2248) );
  inv U1987 ( .in(requested_floor[3]), .out(n2249) );
  inv U1988 ( .in(n2250), .out(\ne_47/AEQB [3]) );
  inv U1989 ( .in(final_floor_elevator1[2]), .out(n2251) );
  inv U1990 ( .in(requested_floor[2]), .out(n2252) );
  inv U1991 ( .in(n2253), .out(\ne_47/AEQB [2]) );
  inv U1992 ( .in(final_floor_elevator1[1]), .out(n2254) );
  inv U1993 ( .in(requested_floor[1]), .out(n2255) );
  inv U1994 ( .in(n2256), .out(\ne_47/AEQB [1]) );
  inv U1995 ( .in(\ne_47/SA ), .out(n2257) );
  inv U1996 ( .in(\ne_47/SB ), .out(n2258) );
  inv U1997 ( .in(n2259), .out(\ne_47/AEQB [63]) );
  inv U1998 ( .in(n2260), .out(\ne_47/LTV [1]) );
  inv U1999 ( .in(final_floor_elevator1[0]), .out(n2261) );
  inv U2000 ( .in(n2262), .out(\ne_47/GTV [1]) );
  inv U2001 ( .in(requested_floor[0]), .out(n2263) );
  inv U2002 ( .in(current_floor_output_elevator2[62]), .out(n2264) );
  inv U2003 ( .in(destination_floor_elevator2[62]), .out(n2265) );
  inv U2004 ( .in(n2266), .out(\eq_47_3/AEQB [62]) );
  inv U2005 ( .in(current_floor_output_elevator2[61]), .out(n2267) );
  inv U2006 ( .in(destination_floor_elevator2[61]), .out(n2268) );
  inv U2007 ( .in(n2269), .out(\eq_47_3/AEQB [61]) );
  inv U2008 ( .in(current_floor_output_elevator2[60]), .out(n2270) );
  inv U2009 ( .in(destination_floor_elevator2[60]), .out(n2271) );
  inv U2010 ( .in(n2272), .out(\eq_47_3/AEQB [60]) );
  inv U2011 ( .in(current_floor_output_elevator2[59]), .out(n2273) );
  inv U2012 ( .in(destination_floor_elevator2[59]), .out(n2274) );
  inv U2013 ( .in(n2275), .out(\eq_47_3/AEQB [59]) );
  inv U2014 ( .in(current_floor_output_elevator2[58]), .out(n2276) );
  inv U2015 ( .in(destination_floor_elevator2[58]), .out(n2277) );
  inv U2016 ( .in(n2278), .out(\eq_47_3/AEQB [58]) );
  inv U2017 ( .in(current_floor_output_elevator2[57]), .out(n2279) );
  inv U2018 ( .in(destination_floor_elevator2[57]), .out(n2280) );
  inv U2019 ( .in(n2281), .out(\eq_47_3/AEQB [57]) );
  inv U2020 ( .in(current_floor_output_elevator2[56]), .out(n2282) );
  inv U2021 ( .in(destination_floor_elevator2[56]), .out(n2283) );
  inv U2022 ( .in(n2284), .out(\eq_47_3/AEQB [56]) );
  inv U2023 ( .in(current_floor_output_elevator2[55]), .out(n2285) );
  inv U2024 ( .in(destination_floor_elevator2[55]), .out(n2286) );
  inv U2025 ( .in(n2287), .out(\eq_47_3/AEQB [55]) );
  inv U2026 ( .in(current_floor_output_elevator2[54]), .out(n2288) );
  inv U2027 ( .in(destination_floor_elevator2[54]), .out(n2289) );
  inv U2028 ( .in(n2290), .out(\eq_47_3/AEQB [54]) );
  inv U2029 ( .in(current_floor_output_elevator2[53]), .out(n2291) );
  inv U2030 ( .in(destination_floor_elevator2[53]), .out(n2292) );
  inv U2031 ( .in(n2293), .out(\eq_47_3/AEQB [53]) );
  inv U2032 ( .in(current_floor_output_elevator2[52]), .out(n2294) );
  inv U2033 ( .in(destination_floor_elevator2[52]), .out(n2295) );
  inv U2034 ( .in(n2296), .out(\eq_47_3/AEQB [52]) );
  inv U2035 ( .in(current_floor_output_elevator2[51]), .out(n2297) );
  inv U2036 ( .in(destination_floor_elevator2[51]), .out(n2298) );
  inv U2037 ( .in(n2299), .out(\eq_47_3/AEQB [51]) );
  inv U2038 ( .in(current_floor_output_elevator2[50]), .out(n2300) );
  inv U2039 ( .in(destination_floor_elevator2[50]), .out(n2301) );
  inv U2040 ( .in(n2302), .out(\eq_47_3/AEQB [50]) );
  inv U2041 ( .in(current_floor_output_elevator2[49]), .out(n2303) );
  inv U2042 ( .in(destination_floor_elevator2[49]), .out(n2304) );
  inv U2043 ( .in(n2305), .out(\eq_47_3/AEQB [49]) );
  inv U2044 ( .in(current_floor_output_elevator2[48]), .out(n2306) );
  inv U2045 ( .in(destination_floor_elevator2[48]), .out(n2307) );
  inv U2046 ( .in(n2308), .out(\eq_47_3/AEQB [48]) );
  inv U2047 ( .in(current_floor_output_elevator2[47]), .out(n2309) );
  inv U2048 ( .in(destination_floor_elevator2[47]), .out(n2310) );
  inv U2049 ( .in(n2311), .out(\eq_47_3/AEQB [47]) );
  inv U2050 ( .in(current_floor_output_elevator2[46]), .out(n2312) );
  inv U2051 ( .in(destination_floor_elevator2[46]), .out(n2313) );
  inv U2052 ( .in(n2314), .out(\eq_47_3/AEQB [46]) );
  inv U2053 ( .in(current_floor_output_elevator2[45]), .out(n2315) );
  inv U2054 ( .in(destination_floor_elevator2[45]), .out(n2316) );
  inv U2055 ( .in(n2317), .out(\eq_47_3/AEQB [45]) );
  inv U2056 ( .in(current_floor_output_elevator2[44]), .out(n2318) );
  inv U2057 ( .in(destination_floor_elevator2[44]), .out(n2319) );
  inv U2058 ( .in(n2320), .out(\eq_47_3/AEQB [44]) );
  inv U2059 ( .in(current_floor_output_elevator2[43]), .out(n2321) );
  inv U2060 ( .in(destination_floor_elevator2[43]), .out(n2322) );
  inv U2061 ( .in(n2323), .out(\eq_47_3/AEQB [43]) );
  inv U2062 ( .in(current_floor_output_elevator2[42]), .out(n2324) );
  inv U2063 ( .in(destination_floor_elevator2[42]), .out(n2325) );
  inv U2064 ( .in(n2326), .out(\eq_47_3/AEQB [42]) );
  inv U2065 ( .in(current_floor_output_elevator2[41]), .out(n2327) );
  inv U2066 ( .in(destination_floor_elevator2[41]), .out(n2328) );
  inv U2067 ( .in(n2329), .out(\eq_47_3/AEQB [41]) );
  inv U2068 ( .in(current_floor_output_elevator2[40]), .out(n2330) );
  inv U2069 ( .in(destination_floor_elevator2[40]), .out(n2331) );
  inv U2070 ( .in(n2332), .out(\eq_47_3/AEQB [40]) );
  inv U2071 ( .in(current_floor_output_elevator2[39]), .out(n2333) );
  inv U2072 ( .in(destination_floor_elevator2[39]), .out(n2334) );
  inv U2073 ( .in(n2335), .out(\eq_47_3/AEQB [39]) );
  inv U2074 ( .in(current_floor_output_elevator2[38]), .out(n2336) );
  inv U2075 ( .in(destination_floor_elevator2[38]), .out(n2337) );
  inv U2076 ( .in(n2338), .out(\eq_47_3/AEQB [38]) );
  inv U2077 ( .in(current_floor_output_elevator2[37]), .out(n2339) );
  inv U2078 ( .in(destination_floor_elevator2[37]), .out(n2340) );
  inv U2079 ( .in(n2341), .out(\eq_47_3/AEQB [37]) );
  inv U2080 ( .in(current_floor_output_elevator2[36]), .out(n2342) );
  inv U2081 ( .in(destination_floor_elevator2[36]), .out(n2343) );
  inv U2082 ( .in(n2344), .out(\eq_47_3/AEQB [36]) );
  inv U2083 ( .in(current_floor_output_elevator2[35]), .out(n2345) );
  inv U2084 ( .in(destination_floor_elevator2[35]), .out(n2346) );
  inv U2085 ( .in(n2347), .out(\eq_47_3/AEQB [35]) );
  inv U2086 ( .in(current_floor_output_elevator2[34]), .out(n2348) );
  inv U2087 ( .in(destination_floor_elevator2[34]), .out(n2349) );
  inv U2088 ( .in(n2350), .out(\eq_47_3/AEQB [34]) );
  inv U2089 ( .in(current_floor_output_elevator2[33]), .out(n2351) );
  inv U2090 ( .in(destination_floor_elevator2[33]), .out(n2352) );
  inv U2091 ( .in(n2353), .out(\eq_47_3/AEQB [33]) );
  inv U2092 ( .in(current_floor_output_elevator2[32]), .out(n2354) );
  inv U2093 ( .in(destination_floor_elevator2[32]), .out(n2355) );
  inv U2094 ( .in(n2356), .out(\eq_47_3/AEQB [32]) );
  inv U2095 ( .in(current_floor_output_elevator2[31]), .out(n2357) );
  inv U2096 ( .in(destination_floor_elevator2[31]), .out(n2358) );
  inv U2097 ( .in(n2359), .out(\eq_47_3/AEQB [31]) );
  inv U2098 ( .in(current_floor_output_elevator2[30]), .out(n2360) );
  inv U2099 ( .in(destination_floor_elevator2[30]), .out(n2361) );
  inv U2100 ( .in(n2362), .out(\eq_47_3/AEQB [30]) );
  inv U2101 ( .in(current_floor_output_elevator2[29]), .out(n2363) );
  inv U2102 ( .in(destination_floor_elevator2[29]), .out(n2364) );
  inv U2103 ( .in(n2365), .out(\eq_47_3/AEQB [29]) );
  inv U2104 ( .in(current_floor_output_elevator2[28]), .out(n2366) );
  inv U2105 ( .in(destination_floor_elevator2[28]), .out(n2367) );
  inv U2106 ( .in(n2368), .out(\eq_47_3/AEQB [28]) );
  inv U2107 ( .in(current_floor_output_elevator2[27]), .out(n2369) );
  inv U2108 ( .in(destination_floor_elevator2[27]), .out(n2370) );
  inv U2109 ( .in(n2371), .out(\eq_47_3/AEQB [27]) );
  inv U2110 ( .in(current_floor_output_elevator2[26]), .out(n2372) );
  inv U2111 ( .in(destination_floor_elevator2[26]), .out(n2373) );
  inv U2112 ( .in(n2374), .out(\eq_47_3/AEQB [26]) );
  inv U2113 ( .in(current_floor_output_elevator2[25]), .out(n2375) );
  inv U2114 ( .in(destination_floor_elevator2[25]), .out(n2376) );
  inv U2115 ( .in(n2377), .out(\eq_47_3/AEQB [25]) );
  inv U2116 ( .in(current_floor_output_elevator2[24]), .out(n2378) );
  inv U2117 ( .in(destination_floor_elevator2[24]), .out(n2379) );
  inv U2118 ( .in(n2380), .out(\eq_47_3/AEQB [24]) );
  inv U2119 ( .in(current_floor_output_elevator2[23]), .out(n2381) );
  inv U2120 ( .in(destination_floor_elevator2[23]), .out(n2382) );
  inv U2121 ( .in(n2383), .out(\eq_47_3/AEQB [23]) );
  inv U2122 ( .in(current_floor_output_elevator2[22]), .out(n2384) );
  inv U2123 ( .in(destination_floor_elevator2[22]), .out(n2385) );
  inv U2124 ( .in(n2386), .out(\eq_47_3/AEQB [22]) );
  inv U2125 ( .in(current_floor_output_elevator2[21]), .out(n2387) );
  inv U2126 ( .in(destination_floor_elevator2[21]), .out(n2388) );
  inv U2127 ( .in(n2389), .out(\eq_47_3/AEQB [21]) );
  inv U2128 ( .in(current_floor_output_elevator2[20]), .out(n2390) );
  inv U2129 ( .in(destination_floor_elevator2[20]), .out(n2391) );
  inv U2130 ( .in(n2392), .out(\eq_47_3/AEQB [20]) );
  inv U2131 ( .in(current_floor_output_elevator2[19]), .out(n2393) );
  inv U2132 ( .in(destination_floor_elevator2[19]), .out(n2394) );
  inv U2133 ( .in(n2395), .out(\eq_47_3/AEQB [19]) );
  inv U2134 ( .in(current_floor_output_elevator2[18]), .out(n2396) );
  inv U2135 ( .in(destination_floor_elevator2[18]), .out(n2397) );
  inv U2136 ( .in(n2398), .out(\eq_47_3/AEQB [18]) );
  inv U2137 ( .in(current_floor_output_elevator2[17]), .out(n2399) );
  inv U2138 ( .in(destination_floor_elevator2[17]), .out(n2400) );
  inv U2139 ( .in(n2401), .out(\eq_47_3/AEQB [17]) );
  inv U2140 ( .in(current_floor_output_elevator2[16]), .out(n2402) );
  inv U2141 ( .in(destination_floor_elevator2[16]), .out(n2403) );
  inv U2142 ( .in(n2404), .out(\eq_47_3/AEQB [16]) );
  inv U2143 ( .in(current_floor_output_elevator2[15]), .out(n2405) );
  inv U2144 ( .in(destination_floor_elevator2[15]), .out(n2406) );
  inv U2145 ( .in(n2407), .out(\eq_47_3/AEQB [15]) );
  inv U2146 ( .in(current_floor_output_elevator2[14]), .out(n2408) );
  inv U2147 ( .in(destination_floor_elevator2[14]), .out(n2409) );
  inv U2148 ( .in(n2410), .out(\eq_47_3/AEQB [14]) );
  inv U2149 ( .in(current_floor_output_elevator2[13]), .out(n2411) );
  inv U2150 ( .in(destination_floor_elevator2[13]), .out(n2412) );
  inv U2151 ( .in(n2413), .out(\eq_47_3/AEQB [13]) );
  inv U2152 ( .in(current_floor_output_elevator2[12]), .out(n2414) );
  inv U2153 ( .in(destination_floor_elevator2[12]), .out(n2415) );
  inv U2154 ( .in(n2416), .out(\eq_47_3/AEQB [12]) );
  inv U2155 ( .in(current_floor_output_elevator2[11]), .out(n2417) );
  inv U2156 ( .in(destination_floor_elevator2[11]), .out(n2418) );
  inv U2157 ( .in(n2419), .out(\eq_47_3/AEQB [11]) );
  inv U2158 ( .in(current_floor_output_elevator2[10]), .out(n2420) );
  inv U2159 ( .in(destination_floor_elevator2[10]), .out(n2421) );
  inv U2160 ( .in(n2422), .out(\eq_47_3/AEQB [10]) );
  inv U2161 ( .in(current_floor_output_elevator2[9]), .out(n2423) );
  inv U2162 ( .in(destination_floor_elevator2[9]), .out(n2424) );
  inv U2163 ( .in(n2425), .out(\eq_47_3/AEQB [9]) );
  inv U2164 ( .in(current_floor_output_elevator2[8]), .out(n2426) );
  inv U2165 ( .in(destination_floor_elevator2[8]), .out(n2427) );
  inv U2166 ( .in(n2428), .out(\eq_47_3/AEQB [8]) );
  inv U2167 ( .in(current_floor_output_elevator2[7]), .out(n2429) );
  inv U2168 ( .in(destination_floor_elevator2[7]), .out(n2430) );
  inv U2169 ( .in(n2431), .out(\eq_47_3/AEQB [7]) );
  inv U2170 ( .in(current_floor_output_elevator2[6]), .out(n2432) );
  inv U2171 ( .in(destination_floor_elevator2[6]), .out(n2433) );
  inv U2172 ( .in(n2434), .out(\eq_47_3/AEQB [6]) );
  inv U2173 ( .in(current_floor_output_elevator2[5]), .out(n2435) );
  inv U2174 ( .in(destination_floor_elevator2[5]), .out(n2436) );
  inv U2175 ( .in(n2437), .out(\eq_47_3/AEQB [5]) );
  inv U2176 ( .in(current_floor_output_elevator2[4]), .out(n2438) );
  inv U2177 ( .in(destination_floor_elevator2[4]), .out(n2439) );
  inv U2178 ( .in(n2440), .out(\eq_47_3/AEQB [4]) );
  inv U2179 ( .in(current_floor_output_elevator2[3]), .out(n2441) );
  inv U2180 ( .in(destination_floor_elevator2[3]), .out(n2442) );
  inv U2181 ( .in(n2443), .out(\eq_47_3/AEQB [3]) );
  inv U2182 ( .in(current_floor_output_elevator2[2]), .out(n2444) );
  inv U2183 ( .in(destination_floor_elevator2[2]), .out(n2445) );
  inv U2184 ( .in(n2446), .out(\eq_47_3/AEQB [2]) );
  inv U2185 ( .in(current_floor_output_elevator2[1]), .out(n2447) );
  inv U2186 ( .in(destination_floor_elevator2[1]), .out(n2448) );
  inv U2187 ( .in(n2449), .out(\eq_47_3/AEQB [1]) );
  inv U2188 ( .in(\eq_47_3/SA ), .out(n2450) );
  inv U2189 ( .in(\eq_47_3/SB ), .out(n2451) );
  inv U2190 ( .in(n2452), .out(\eq_47_3/AEQB [63]) );
  inv U2191 ( .in(n2453), .out(\eq_47_3/LTV [1]) );
  inv U2192 ( .in(current_floor_output_elevator2[0]), .out(n2454) );
  inv U2193 ( .in(n2455), .out(\eq_47_3/GTV [1]) );
  inv U2194 ( .in(destination_floor_elevator2[0]), .out(n2456) );
  inv U2195 ( .in(N156), .out(n2457) );
  inv U2196 ( .in(N92), .out(n2458) );
  inv U2197 ( .in(n2459), .out(\r125/AEQB [62]) );
  inv U2198 ( .in(N157), .out(n2460) );
  inv U2199 ( .in(N93), .out(n2461) );
  inv U2200 ( .in(n2462), .out(\r125/AEQB [61]) );
  inv U2201 ( .in(N158), .out(n2463) );
  inv U2202 ( .in(N94), .out(n2464) );
  inv U2203 ( .in(n2465), .out(\r125/AEQB [60]) );
  inv U2204 ( .in(N159), .out(n2466) );
  inv U2205 ( .in(N95), .out(n2467) );
  inv U2206 ( .in(n2468), .out(\r125/AEQB [59]) );
  inv U2207 ( .in(N160), .out(n2469) );
  inv U2208 ( .in(N96), .out(n2470) );
  inv U2209 ( .in(n2471), .out(\r125/AEQB [58]) );
  inv U2210 ( .in(N161), .out(n2472) );
  inv U2211 ( .in(N97), .out(n2473) );
  inv U2212 ( .in(n2474), .out(\r125/AEQB [57]) );
  inv U2213 ( .in(N162), .out(n2475) );
  inv U2214 ( .in(N98), .out(n2476) );
  inv U2215 ( .in(n2477), .out(\r125/AEQB [56]) );
  inv U2216 ( .in(N163), .out(n2478) );
  inv U2217 ( .in(N99), .out(n2479) );
  inv U2218 ( .in(n2480), .out(\r125/AEQB [55]) );
  inv U2219 ( .in(N164), .out(n2481) );
  inv U2220 ( .in(N100), .out(n2482) );
  inv U2221 ( .in(n2483), .out(\r125/AEQB [54]) );
  inv U2222 ( .in(N165), .out(n2484) );
  inv U2223 ( .in(N101), .out(n2485) );
  inv U2224 ( .in(n2486), .out(\r125/AEQB [53]) );
  inv U2225 ( .in(N166), .out(n2487) );
  inv U2226 ( .in(N102), .out(n2488) );
  inv U2227 ( .in(n2489), .out(\r125/AEQB [52]) );
  inv U2228 ( .in(N167), .out(n2490) );
  inv U2229 ( .in(N103), .out(n2491) );
  inv U2230 ( .in(n2492), .out(\r125/AEQB [51]) );
  inv U2231 ( .in(N168), .out(n2493) );
  inv U2232 ( .in(N104), .out(n2494) );
  inv U2233 ( .in(n2495), .out(\r125/AEQB [50]) );
  inv U2234 ( .in(N169), .out(n2496) );
  inv U2235 ( .in(N105), .out(n2497) );
  inv U2236 ( .in(n2498), .out(\r125/AEQB [49]) );
  inv U2237 ( .in(N170), .out(n2499) );
  inv U2238 ( .in(N106), .out(n2500) );
  inv U2239 ( .in(n2501), .out(\r125/AEQB [48]) );
  inv U2240 ( .in(N171), .out(n2502) );
  inv U2241 ( .in(N107), .out(n2503) );
  inv U2242 ( .in(n2504), .out(\r125/AEQB [47]) );
  inv U2243 ( .in(N172), .out(n2505) );
  inv U2244 ( .in(N108), .out(n2506) );
  inv U2245 ( .in(n2507), .out(\r125/AEQB [46]) );
  inv U2246 ( .in(N173), .out(n2508) );
  inv U2247 ( .in(N109), .out(n2509) );
  inv U2248 ( .in(n2510), .out(\r125/AEQB [45]) );
  inv U2249 ( .in(N174), .out(n2511) );
  inv U2250 ( .in(N110), .out(n2512) );
  inv U2251 ( .in(n2513), .out(\r125/AEQB [44]) );
  inv U2252 ( .in(N175), .out(n2514) );
  inv U2253 ( .in(N111), .out(n2515) );
  inv U2254 ( .in(n2516), .out(\r125/AEQB [43]) );
  inv U2255 ( .in(N176), .out(n2517) );
  inv U2256 ( .in(N112), .out(n2518) );
  inv U2257 ( .in(n2519), .out(\r125/AEQB [42]) );
  inv U2258 ( .in(N177), .out(n2520) );
  inv U2259 ( .in(N113), .out(n2521) );
  inv U2260 ( .in(n2522), .out(\r125/AEQB [41]) );
  inv U2261 ( .in(N178), .out(n2523) );
  inv U2262 ( .in(N114), .out(n2524) );
  inv U2263 ( .in(n2525), .out(\r125/AEQB [40]) );
  inv U2264 ( .in(N179), .out(n2526) );
  inv U2265 ( .in(N115), .out(n2527) );
  inv U2266 ( .in(n2528), .out(\r125/AEQB [39]) );
  inv U2267 ( .in(N180), .out(n2529) );
  inv U2268 ( .in(N116), .out(n2530) );
  inv U2269 ( .in(n2531), .out(\r125/AEQB [38]) );
  inv U2270 ( .in(N181), .out(n2532) );
  inv U2271 ( .in(N117), .out(n2533) );
  inv U2272 ( .in(n2534), .out(\r125/AEQB [37]) );
  inv U2273 ( .in(N182), .out(n2535) );
  inv U2274 ( .in(N118), .out(n2536) );
  inv U2275 ( .in(n2537), .out(\r125/AEQB [36]) );
  inv U2276 ( .in(N183), .out(n2538) );
  inv U2277 ( .in(N119), .out(n2539) );
  inv U2278 ( .in(n2540), .out(\r125/AEQB [35]) );
  inv U2279 ( .in(N184), .out(n2541) );
  inv U2280 ( .in(N120), .out(n2542) );
  inv U2281 ( .in(n2543), .out(\r125/AEQB [34]) );
  inv U2282 ( .in(N185), .out(n2544) );
  inv U2283 ( .in(N121), .out(n2545) );
  inv U2284 ( .in(n2546), .out(\r125/AEQB [33]) );
  inv U2285 ( .in(N186), .out(n2547) );
  inv U2286 ( .in(N122), .out(n2548) );
  inv U2287 ( .in(n2549), .out(\r125/AEQB [32]) );
  inv U2288 ( .in(N187), .out(n2550) );
  inv U2289 ( .in(N123), .out(n2551) );
  inv U2290 ( .in(n2552), .out(\r125/AEQB [31]) );
  inv U2291 ( .in(N188), .out(n2553) );
  inv U2292 ( .in(N124), .out(n2554) );
  inv U2293 ( .in(n2555), .out(\r125/AEQB [30]) );
  inv U2294 ( .in(N189), .out(n2556) );
  inv U2295 ( .in(N125), .out(n2557) );
  inv U2296 ( .in(n2558), .out(\r125/AEQB [29]) );
  inv U2297 ( .in(N190), .out(n2559) );
  inv U2298 ( .in(N126), .out(n2560) );
  inv U2299 ( .in(n2561), .out(\r125/AEQB [28]) );
  inv U2300 ( .in(N191), .out(n2562) );
  inv U2301 ( .in(N127), .out(n2563) );
  inv U2302 ( .in(n2564), .out(\r125/AEQB [27]) );
  inv U2303 ( .in(N192), .out(n2565) );
  inv U2304 ( .in(N128), .out(n2566) );
  inv U2305 ( .in(n2567), .out(\r125/AEQB [26]) );
  inv U2306 ( .in(N193), .out(n2568) );
  inv U2307 ( .in(N129), .out(n2569) );
  inv U2308 ( .in(n2570), .out(\r125/AEQB [25]) );
  inv U2309 ( .in(N194), .out(n2571) );
  inv U2310 ( .in(N130), .out(n2572) );
  inv U2311 ( .in(n2573), .out(\r125/AEQB [24]) );
  inv U2312 ( .in(N195), .out(n2574) );
  inv U2313 ( .in(N131), .out(n2575) );
  inv U2314 ( .in(n2576), .out(\r125/AEQB [23]) );
  inv U2315 ( .in(N196), .out(n2577) );
  inv U2316 ( .in(N132), .out(n2578) );
  inv U2317 ( .in(n2579), .out(\r125/AEQB [22]) );
  inv U2318 ( .in(N197), .out(n2580) );
  inv U2319 ( .in(N133), .out(n2581) );
  inv U2320 ( .in(n2582), .out(\r125/AEQB [21]) );
  inv U2321 ( .in(N198), .out(n2583) );
  inv U2322 ( .in(N134), .out(n2584) );
  inv U2323 ( .in(n2585), .out(\r125/AEQB [20]) );
  inv U2324 ( .in(N199), .out(n2586) );
  inv U2325 ( .in(N135), .out(n2587) );
  inv U2326 ( .in(n2588), .out(\r125/AEQB [19]) );
  inv U2327 ( .in(N200), .out(n2589) );
  inv U2328 ( .in(N136), .out(n2590) );
  inv U2329 ( .in(n2591), .out(\r125/AEQB [18]) );
  inv U2330 ( .in(N201), .out(n2592) );
  inv U2331 ( .in(N137), .out(n2593) );
  inv U2332 ( .in(n2594), .out(\r125/AEQB [17]) );
  inv U2333 ( .in(N202), .out(n2595) );
  inv U2334 ( .in(N138), .out(n2596) );
  inv U2335 ( .in(n2597), .out(\r125/AEQB [16]) );
  inv U2336 ( .in(N203), .out(n2598) );
  inv U2337 ( .in(N139), .out(n2599) );
  inv U2338 ( .in(n2600), .out(\r125/AEQB [15]) );
  inv U2339 ( .in(N204), .out(n2601) );
  inv U2340 ( .in(N140), .out(n2602) );
  inv U2341 ( .in(n2603), .out(\r125/AEQB [14]) );
  inv U2342 ( .in(N205), .out(n2604) );
  inv U2343 ( .in(N141), .out(n2605) );
  inv U2344 ( .in(n2606), .out(\r125/AEQB [13]) );
  inv U2345 ( .in(N206), .out(n2607) );
  inv U2346 ( .in(N142), .out(n2608) );
  inv U2347 ( .in(n2609), .out(\r125/AEQB [12]) );
  inv U2348 ( .in(N207), .out(n2610) );
  inv U2349 ( .in(N143), .out(n2611) );
  inv U2350 ( .in(n2612), .out(\r125/AEQB [11]) );
  inv U2351 ( .in(N208), .out(n2613) );
  inv U2352 ( .in(N144), .out(n2614) );
  inv U2353 ( .in(n2615), .out(\r125/AEQB [10]) );
  inv U2354 ( .in(N209), .out(n2616) );
  inv U2355 ( .in(N145), .out(n2617) );
  inv U2356 ( .in(n2618), .out(\r125/AEQB [9]) );
  inv U2357 ( .in(N210), .out(n2619) );
  inv U2358 ( .in(N146), .out(n2620) );
  inv U2359 ( .in(n2621), .out(\r125/AEQB [8]) );
  inv U2360 ( .in(N211), .out(n2622) );
  inv U2361 ( .in(N147), .out(n2623) );
  inv U2362 ( .in(n2624), .out(\r125/AEQB [7]) );
  inv U2363 ( .in(N212), .out(n2625) );
  inv U2364 ( .in(N148), .out(n2626) );
  inv U2365 ( .in(n2627), .out(\r125/AEQB [6]) );
  inv U2366 ( .in(N213), .out(n2628) );
  inv U2367 ( .in(N149), .out(n2629) );
  inv U2368 ( .in(n2630), .out(\r125/AEQB [5]) );
  inv U2369 ( .in(N214), .out(n2631) );
  inv U2370 ( .in(N150), .out(n2632) );
  inv U2371 ( .in(n2633), .out(\r125/AEQB [4]) );
  inv U2372 ( .in(N215), .out(n2634) );
  inv U2373 ( .in(N151), .out(n2635) );
  inv U2374 ( .in(n2636), .out(\r125/AEQB [3]) );
  inv U2375 ( .in(N216), .out(n2637) );
  inv U2376 ( .in(N152), .out(n2638) );
  inv U2377 ( .in(n2639), .out(\r125/AEQB [2]) );
  inv U2378 ( .in(N217), .out(n2640) );
  inv U2379 ( .in(N153), .out(n2641) );
  inv U2380 ( .in(n2642), .out(\r125/AEQB [1]) );
  inv U2381 ( .in(\r125/SA ), .out(n2643) );
  inv U2382 ( .in(\r125/SB ), .out(n2644) );
  inv U2383 ( .in(n2645), .out(\r125/AEQB [63]) );
  inv U2384 ( .in(n2646), .out(\r125/LTV [1]) );
  inv U2385 ( .in(N218), .out(n2647) );
  inv U2386 ( .in(n2648), .out(\r125/GTV [1]) );
  inv U2387 ( .in(N154), .out(n2649) );
  inv U2388 ( .in(N440), .out(n2650) );
  inv U2389 ( .in(N376), .out(n2651) );
  inv U2390 ( .in(n2652), .out(\r126/AEQB [62]) );
  inv U2391 ( .in(N441), .out(n2653) );
  inv U2392 ( .in(N377), .out(n2654) );
  inv U2393 ( .in(n2655), .out(\r126/AEQB [61]) );
  inv U2394 ( .in(N442), .out(n2656) );
  inv U2395 ( .in(N378), .out(n2657) );
  inv U2396 ( .in(n2658), .out(\r126/AEQB [60]) );
  inv U2397 ( .in(N443), .out(n2659) );
  inv U2398 ( .in(N379), .out(n2660) );
  inv U2399 ( .in(n2661), .out(\r126/AEQB [59]) );
  inv U2400 ( .in(N444), .out(n2662) );
  inv U2401 ( .in(N380), .out(n2663) );
  inv U2402 ( .in(n2664), .out(\r126/AEQB [58]) );
  inv U2403 ( .in(N445), .out(n2665) );
  inv U2404 ( .in(N381), .out(n2666) );
  inv U2405 ( .in(n2667), .out(\r126/AEQB [57]) );
  inv U2406 ( .in(N446), .out(n2668) );
  inv U2407 ( .in(N382), .out(n2669) );
  inv U2408 ( .in(n2670), .out(\r126/AEQB [56]) );
  inv U2409 ( .in(N447), .out(n2671) );
  inv U2410 ( .in(N383), .out(n2672) );
  inv U2411 ( .in(n2673), .out(\r126/AEQB [55]) );
  inv U2412 ( .in(N448), .out(n2674) );
  inv U2413 ( .in(N384), .out(n2675) );
  inv U2414 ( .in(n2676), .out(\r126/AEQB [54]) );
  inv U2415 ( .in(N449), .out(n2677) );
  inv U2416 ( .in(N385), .out(n2678) );
  inv U2417 ( .in(n2679), .out(\r126/AEQB [53]) );
  inv U2418 ( .in(N450), .out(n2680) );
  inv U2419 ( .in(N386), .out(n2681) );
  inv U2420 ( .in(n2682), .out(\r126/AEQB [52]) );
  inv U2421 ( .in(N451), .out(n2683) );
  inv U2422 ( .in(N387), .out(n2684) );
  inv U2423 ( .in(n2685), .out(\r126/AEQB [51]) );
  inv U2424 ( .in(N452), .out(n2686) );
  inv U2425 ( .in(N388), .out(n2687) );
  inv U2426 ( .in(n2688), .out(\r126/AEQB [50]) );
  inv U2427 ( .in(N453), .out(n2689) );
  inv U2428 ( .in(N389), .out(n2690) );
  inv U2429 ( .in(n2691), .out(\r126/AEQB [49]) );
  inv U2430 ( .in(N454), .out(n2692) );
  inv U2431 ( .in(N390), .out(n2693) );
  inv U2432 ( .in(n2694), .out(\r126/AEQB [48]) );
  inv U2433 ( .in(N455), .out(n2695) );
  inv U2434 ( .in(N391), .out(n2696) );
  inv U2435 ( .in(n2697), .out(\r126/AEQB [47]) );
  inv U2436 ( .in(N456), .out(n2698) );
  inv U2437 ( .in(N392), .out(n2699) );
  inv U2438 ( .in(n2700), .out(\r126/AEQB [46]) );
  inv U2439 ( .in(N457), .out(n2701) );
  inv U2440 ( .in(N393), .out(n2702) );
  inv U2441 ( .in(n2703), .out(\r126/AEQB [45]) );
  inv U2442 ( .in(N458), .out(n2704) );
  inv U2443 ( .in(N394), .out(n2705) );
  inv U2444 ( .in(n2706), .out(\r126/AEQB [44]) );
  inv U2445 ( .in(N459), .out(n2707) );
  inv U2446 ( .in(N395), .out(n2708) );
  inv U2447 ( .in(n2709), .out(\r126/AEQB [43]) );
  inv U2448 ( .in(N460), .out(n2710) );
  inv U2449 ( .in(N396), .out(n2711) );
  inv U2450 ( .in(n2712), .out(\r126/AEQB [42]) );
  inv U2451 ( .in(N461), .out(n2713) );
  inv U2452 ( .in(N397), .out(n2714) );
  inv U2453 ( .in(n2715), .out(\r126/AEQB [41]) );
  inv U2454 ( .in(N462), .out(n2716) );
  inv U2455 ( .in(N398), .out(n2717) );
  inv U2456 ( .in(n2718), .out(\r126/AEQB [40]) );
  inv U2457 ( .in(N463), .out(n2719) );
  inv U2458 ( .in(N399), .out(n2720) );
  inv U2459 ( .in(n2721), .out(\r126/AEQB [39]) );
  inv U2460 ( .in(N464), .out(n2722) );
  inv U2461 ( .in(N400), .out(n2723) );
  inv U2462 ( .in(n2724), .out(\r126/AEQB [38]) );
  inv U2463 ( .in(N465), .out(n2725) );
  inv U2464 ( .in(N401), .out(n2726) );
  inv U2465 ( .in(n2727), .out(\r126/AEQB [37]) );
  inv U2466 ( .in(N466), .out(n2728) );
  inv U2467 ( .in(N402), .out(n2729) );
  inv U2468 ( .in(n2730), .out(\r126/AEQB [36]) );
  inv U2469 ( .in(N467), .out(n2731) );
  inv U2470 ( .in(N403), .out(n2732) );
  inv U2471 ( .in(n2733), .out(\r126/AEQB [35]) );
  inv U2472 ( .in(N468), .out(n2734) );
  inv U2473 ( .in(N404), .out(n2735) );
  inv U2474 ( .in(n2736), .out(\r126/AEQB [34]) );
  inv U2475 ( .in(N469), .out(n2737) );
  inv U2476 ( .in(N405), .out(n2738) );
  inv U2477 ( .in(n2739), .out(\r126/AEQB [33]) );
  inv U2478 ( .in(N470), .out(n2740) );
  inv U2479 ( .in(N406), .out(n2741) );
  inv U2480 ( .in(n2742), .out(\r126/AEQB [32]) );
  inv U2481 ( .in(N471), .out(n2743) );
  inv U2482 ( .in(N407), .out(n2744) );
  inv U2483 ( .in(n2745), .out(\r126/AEQB [31]) );
  inv U2484 ( .in(N472), .out(n2746) );
  inv U2485 ( .in(N408), .out(n2747) );
  inv U2486 ( .in(n2748), .out(\r126/AEQB [30]) );
  inv U2487 ( .in(N473), .out(n2749) );
  inv U2488 ( .in(N409), .out(n2750) );
  inv U2489 ( .in(n2751), .out(\r126/AEQB [29]) );
  inv U2490 ( .in(N474), .out(n2752) );
  inv U2491 ( .in(N410), .out(n2753) );
  inv U2492 ( .in(n2754), .out(\r126/AEQB [28]) );
  inv U2493 ( .in(N475), .out(n2755) );
  inv U2494 ( .in(N411), .out(n2756) );
  inv U2495 ( .in(n2757), .out(\r126/AEQB [27]) );
  inv U2496 ( .in(N476), .out(n2758) );
  inv U2497 ( .in(N412), .out(n2759) );
  inv U2498 ( .in(n2760), .out(\r126/AEQB [26]) );
  inv U2499 ( .in(N477), .out(n2761) );
  inv U2500 ( .in(N413), .out(n2762) );
  inv U2501 ( .in(n2763), .out(\r126/AEQB [25]) );
  inv U2502 ( .in(N478), .out(n2764) );
  inv U2503 ( .in(N414), .out(n2765) );
  inv U2504 ( .in(n2766), .out(\r126/AEQB [24]) );
  inv U2505 ( .in(N479), .out(n2767) );
  inv U2506 ( .in(N415), .out(n2768) );
  inv U2507 ( .in(n2769), .out(\r126/AEQB [23]) );
  inv U2508 ( .in(N480), .out(n2770) );
  inv U2509 ( .in(N416), .out(n2771) );
  inv U2510 ( .in(n2772), .out(\r126/AEQB [22]) );
  inv U2511 ( .in(N481), .out(n2773) );
  inv U2512 ( .in(N417), .out(n2774) );
  inv U2513 ( .in(n2775), .out(\r126/AEQB [21]) );
  inv U2514 ( .in(N482), .out(n2776) );
  inv U2515 ( .in(N418), .out(n2777) );
  inv U2516 ( .in(n2778), .out(\r126/AEQB [20]) );
  inv U2517 ( .in(N483), .out(n2779) );
  inv U2518 ( .in(N419), .out(n2780) );
  inv U2519 ( .in(n2781), .out(\r126/AEQB [19]) );
  inv U2520 ( .in(N484), .out(n2782) );
  inv U2521 ( .in(N420), .out(n2783) );
  inv U2522 ( .in(n2784), .out(\r126/AEQB [18]) );
  inv U2523 ( .in(N485), .out(n2785) );
  inv U2524 ( .in(N421), .out(n2786) );
  inv U2525 ( .in(n2787), .out(\r126/AEQB [17]) );
  inv U2526 ( .in(N486), .out(n2788) );
  inv U2527 ( .in(N422), .out(n2789) );
  inv U2528 ( .in(n2790), .out(\r126/AEQB [16]) );
  inv U2529 ( .in(N487), .out(n2791) );
  inv U2530 ( .in(N423), .out(n2792) );
  inv U2531 ( .in(n2793), .out(\r126/AEQB [15]) );
  inv U2532 ( .in(N488), .out(n2794) );
  inv U2533 ( .in(N424), .out(n2795) );
  inv U2534 ( .in(n2796), .out(\r126/AEQB [14]) );
  inv U2535 ( .in(N489), .out(n2797) );
  inv U2536 ( .in(N425), .out(n2798) );
  inv U2537 ( .in(n2799), .out(\r126/AEQB [13]) );
  inv U2538 ( .in(N490), .out(n2800) );
  inv U2539 ( .in(N426), .out(n2801) );
  inv U2540 ( .in(n2802), .out(\r126/AEQB [12]) );
  inv U2541 ( .in(N491), .out(n2803) );
  inv U2542 ( .in(N427), .out(n2804) );
  inv U2543 ( .in(n2805), .out(\r126/AEQB [11]) );
  inv U2544 ( .in(N492), .out(n2806) );
  inv U2545 ( .in(N428), .out(n2807) );
  inv U2546 ( .in(n2808), .out(\r126/AEQB [10]) );
  inv U2547 ( .in(N493), .out(n2809) );
  inv U2548 ( .in(N429), .out(n2810) );
  inv U2549 ( .in(n2811), .out(\r126/AEQB [9]) );
  inv U2550 ( .in(N494), .out(n2812) );
  inv U2551 ( .in(N430), .out(n2813) );
  inv U2552 ( .in(n2814), .out(\r126/AEQB [8]) );
  inv U2553 ( .in(N495), .out(n2815) );
  inv U2554 ( .in(N431), .out(n2816) );
  inv U2555 ( .in(n2817), .out(\r126/AEQB [7]) );
  inv U2556 ( .in(N496), .out(n2818) );
  inv U2557 ( .in(N432), .out(n2819) );
  inv U2558 ( .in(n2820), .out(\r126/AEQB [6]) );
  inv U2559 ( .in(N497), .out(n2821) );
  inv U2560 ( .in(N433), .out(n2822) );
  inv U2561 ( .in(n2823), .out(\r126/AEQB [5]) );
  inv U2562 ( .in(N498), .out(n2824) );
  inv U2563 ( .in(N434), .out(n2825) );
  inv U2564 ( .in(n2826), .out(\r126/AEQB [4]) );
  inv U2565 ( .in(N499), .out(n2827) );
  inv U2566 ( .in(N435), .out(n2828) );
  inv U2567 ( .in(n2829), .out(\r126/AEQB [3]) );
  inv U2568 ( .in(N500), .out(n2830) );
  inv U2569 ( .in(N436), .out(n2831) );
  inv U2570 ( .in(n2832), .out(\r126/AEQB [2]) );
  inv U2571 ( .in(N501), .out(n2833) );
  inv U2572 ( .in(N437), .out(n2834) );
  inv U2573 ( .in(n2835), .out(\r126/AEQB [1]) );
  inv U2574 ( .in(\r126/SA ), .out(n2836) );
  inv U2575 ( .in(\r126/SB ), .out(n2837) );
  inv U2576 ( .in(n2838), .out(\r126/AEQB [63]) );
  inv U2577 ( .in(n2839), .out(\r126/LTV [1]) );
  inv U2578 ( .in(N502), .out(n2840) );
  inv U2579 ( .in(n2841), .out(\r126/GTV [1]) );
  inv U2580 ( .in(N438), .out(n2842) );
endmodule

