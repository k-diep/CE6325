* File: xor2.pex.sp
* Created: Fri Oct 27 14:32:42 2023
* Program "Calibre xRC"
* Version "v2013.2_18.13"
* 
.include "xor2.pex.sp.pex"
.subckt xor2  VSS OUT VDD B A
* 
* A	A
* B	B
* VDD	VDD
* OUT	OUT
* VSS	VSS
XD0_noxref N_VSS_D0_noxref_pos N_VDD_D0_noxref_neg DIODENWX  AREA=8.01852e-12
+ PERIM=1.154e-05
XMMN3 N_NET9_MMN3_d N_B_MMN3_g N_VSS_MMN3_s N_VSS_D0_noxref_pos NFET L=6.5e-08
+ W=5.6e-07 AD=1.2964e-13 AS=1.8984e-13 PD=1.023e-06 PS=1.798e-06 NRD=0.282143
+ NRS=0.317857 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=3.39e-07
+ SB=2.283e-06 SD=0 PANW1=7.54e-15 PANW2=3.25e-15 PANW3=3.25e-15 PANW4=3.25e-15
+ PANW5=3.25e-15 PANW6=6.5e-15 PANW7=9.36e-15 PANW8=0 PANW9=0 PANW10=0
XMMN2 N_NET9_MMN3_d N_A_MMN2_g N_VSS_MMN2_s N_VSS_D0_noxref_pos NFET L=6.5e-08
+ W=5.6e-07 AD=1.2964e-13 AS=1.3104e-13 PD=1.023e-06 PS=1.028e-06 NRD=0.544643
+ NRS=0.289286 M=1 NF=1 CNR_SWITCH=1 PCCRIT=0 PAR=1 PTWELL=0 SA=8.67e-07
+ SB=1.755e-06 SD=0 PANW1=7.54e-15 PANW2=3.25e-15 PANW3=3.25e-15 PANW4=3.25e-15
+ PANW5=3.25e-15 PANW6=6.5e-15 PANW7=9.36e-15 PANW8=0 PANW9=0 PANW10=0
XMMN0 N_OUT_MMN0_d N_NET9_MMN0_g N_VSS_MMN2_s N_VSS_D0_noxref_pos NFET
+ L=6.5e-08 W=5.6e-07 AD=1.2992e-13 AS=1.3104e-13 PD=1.024e-06 PS=1.028e-06
+ NRD=0.289286 NRS=0.546429 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0
+ SA=1.4e-06 SB=1.222e-06 SD=0 PANW1=7.54e-15 PANW2=3.25e-15 PANW3=3.25e-15
+ PANW4=3.25e-15 PANW5=3.25e-15 PANW6=6.5e-15 PANW7=9.36e-15 PANW8=0 PANW9=0
+ PANW10=0
XMMN1 N_OUT_MMN0_d N_A_MMN1_g NET26 N_VSS_D0_noxref_pos NFET L=6.5e-08
+ W=5.6e-07 AD=1.2992e-13 AS=1.3076e-13 PD=1.024e-06 PS=1.027e-06 NRD=0.539286
+ NRS=0.416964 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=1.929e-06
+ SB=6.93e-07 SD=0 PANW1=7.54e-15 PANW2=3.25e-15 PANW3=3.25e-15 PANW4=3.25e-15
+ PANW5=3.25e-15 PANW6=6.5e-15 PANW7=9.36e-15 PANW8=0 PANW9=0 PANW10=0
XMMN4 NET26 N_B_MMN4_g N_VSS_MMN4_s N_VSS_D0_noxref_pos NFET L=6.5e-08
+ W=5.6e-07 AD=1.3076e-13 AS=9.016e-14 PD=1.027e-06 PS=1.442e-06 NRD=0.416964
+ NRS=0.178571 M=1 NF=1 CNR_SWITCH=1 PCCRIT=0 PAR=1 PTWELL=0 SA=2.461e-06
+ SB=1.61e-07 SD=0 PANW1=7.54e-15 PANW2=3.25e-15 PANW3=3.25e-15 PANW4=3.25e-15
+ PANW5=3.25e-15 PANW6=6.5e-15 PANW7=9.36e-15 PANW8=0 PANW9=0 PANW10=0
XMMP0 N_NET9_MMP0_d N_B_MMP0_g NET27 N_VDD_D0_noxref_neg PFET L=6.5e-08
+ W=9.6e-07 AD=3.2544e-13 AS=2.2224e-13 PD=2.598e-06 PS=1.423e-06 NRD=0.185417
+ NRS=0.241146 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=3.39e-07
+ SB=2.283e-06 SD=0 PANW1=0 PANW2=0 PANW3=1.885e-15 PANW4=3.25e-15
+ PANW5=3.25e-15 PANW6=6.5e-15 PANW7=7.54e-14 PANW8=1.3e-14 PANW9=4.7385e-14
+ PANW10=3.653e-14
XMMP3 NET27 N_A_MMP3_g N_VDD_MMP3_s N_VDD_D0_noxref_neg PFET L=6.5e-08
+ W=9.6e-07 AD=2.2224e-13 AS=2.2464e-13 PD=1.423e-06 PS=1.428e-06 NRD=0.241146
+ NRS=0.16875 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=8.67e-07
+ SB=1.755e-06 SD=0 PANW1=0 PANW2=0 PANW3=1.885e-15 PANW4=3.25e-15
+ PANW5=3.25e-15 PANW6=6.5e-15 PANW7=1.3e-14 PANW8=1.3e-14 PANW9=1.09785e-13
+ PANW10=3.653e-14
XMMP1 N_NET14_MMP1_d N_NET9_MMP1_g N_VDD_MMP3_s N_VDD_D0_noxref_neg PFET
+ L=6.5e-08 W=9.6e-07 AD=2.2272e-13 AS=2.2464e-13 PD=1.424e-06 PS=1.428e-06
+ NRD=0.16875 NRS=0.31875 M=1 NF=1 CNR_SWITCH=2 PCCRIT=0 PAR=1 PTWELL=1
+ SA=1.4e-06 SB=1.222e-06 SD=0 PANW1=0 PANW2=0 PANW3=1.885e-15 PANW4=3.25e-15
+ PANW5=3.25e-15 PANW6=6.5e-15 PANW7=1.3e-14 PANW8=1.3e-14 PANW9=4.7385e-14
+ PANW10=1.6133e-13
XMMP2 N_OUT_MMP2_d N_A_MMP2_g N_NET14_MMP1_d N_VDD_D0_noxref_neg PFET L=6.5e-08
+ W=9.6e-07 AD=2.2416e-13 AS=2.2272e-13 PD=1.427e-06 PS=1.424e-06 NRD=0.182292
+ NRS=0.314583 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=1.929e-06
+ SB=6.93e-07 SD=0 PANW1=0 PANW2=0 PANW3=1.885e-15 PANW4=3.25e-15 PANW5=3.25e-15
+ PANW6=6.5e-15 PANW7=1.3e-14 PANW8=1.3e-14 PANW9=1.09785e-13 PANW10=3.653e-14
XMMP4 N_OUT_MMP2_d N_B_MMP4_g N_NET14_MMP4_s N_VDD_D0_noxref_neg PFET L=6.5e-08
+ W=9.6e-07 AD=2.2416e-13 AS=1.5456e-13 PD=1.427e-06 PS=2.242e-06 NRD=0.304167
+ NRS=0.105208 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=2.461e-06
+ SB=1.61e-07 SD=0 PANW1=0 PANW2=0 PANW3=1.885e-15 PANW4=3.25e-15 PANW5=3.25e-15
+ PANW6=6.89e-14 PANW7=1.3e-14 PANW8=1.3e-14 PANW9=4.7385e-14 PANW10=3.653e-14
*
.include "xor2.pex.sp.XOR2.pxi"
*
.ends
*
*
