* File: /home/012/k/kt/ktd170030/cad/gf65/NOR3_PEX/nor3.pex.sp
* Created: Thu Oct 26 18:23:13 2023
* Program "Calibre xRC"
* Version "v2013.2_18.13"
* 
.include "/home/012/k/kt/ktd170030/cad/gf65/NOR3_PEX/nor3.pex.sp.pex"
.subckt nor3  VSS OUT VDD A B C
* 
* C	C
* B	B
* A	A
* VDD	VDD
* OUT	OUT
* VSS	VSS
XD0_noxref N_VSS_D0_noxref_pos N_VDD_D0_noxref_neg DIODENWX  AREA=1.04744e-11
+ PERIM=1.3484e-05
XMMN3 N_OUT_MMN3_d N_A_MMN3_g N_VSS_MMN3_s N_VSS_D0_noxref_pos NFET L=6.5e-08
+ W=5.6e-07 AD=1.246e-13 AS=1.3552e-13 PD=1.005e-06 PS=1.604e-06 NRD=0.178571
+ NRS=0.178571 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=2.42e-07
+ SB=1.261e-06 SD=0 PANW1=0 PANW2=0 PANW3=2.34e-15 PANW4=3.25e-15 PANW5=3.25e-15
+ PANW6=6.5e-15 PANW7=1.3e-14 PANW8=8.06e-15 PANW9=0 PANW10=0
XMMN0 N_OUT_MMN3_d N_B_MMN0_g N_VSS_MMN0_s N_VSS_D0_noxref_pos NFET L=6.5e-08
+ W=5.6e-07 AD=1.246e-13 AS=1.274e-13 PD=1.005e-06 PS=1.015e-06 NRD=0.616071
+ NRS=0.414286 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=7.52e-07
+ SB=7.51e-07 SD=0 PANW1=0 PANW2=0 PANW3=2.34e-15 PANW4=3.25e-15 PANW5=3.25e-15
+ PANW6=6.5e-15 PANW7=1.3e-14 PANW8=8.06e-15 PANW9=0 PANW10=0
XMMN2 N_OUT_MMN2_d N_C_MMN2_g N_VSS_MMN0_s N_VSS_D0_noxref_pos NFET L=6.5e-08
+ W=5.6e-07 AD=1.2936e-13 AS=1.274e-13 PD=1.582e-06 PS=1.015e-06 NRD=0.196429
+ NRS=0.398214 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=0 SA=1.272e-06
+ SB=2.31e-07 SD=0 PANW1=0 PANW2=0 PANW3=2.34e-15 PANW4=3.25e-15 PANW5=3.25e-15
+ PANW6=6.5e-15 PANW7=1.3e-14 PANW8=8.06e-15 PANW9=0 PANW10=0
XMMP0 NET16 N_A_MMP0_g N_VDD_MMP0_s N_VDD_D0_noxref_neg PFET L=6.5e-08
+ W=9.6e-07 AD=2.136e-13 AS=2.3232e-13 PD=1.405e-06 PS=2.404e-06 NRD=0.231771
+ NRS=0.104167 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=2.42e-07
+ SB=1.261e-06 SD=0 PANW1=0 PANW2=0 PANW3=1.885e-15 PANW4=3.25e-15
+ PANW5=3.25e-15 PANW6=6.5e-15 PANW7=1.3e-14 PANW8=1.3e-14 PANW9=4.121e-14
+ PANW10=1.014e-13
XMMP1 NET016 N_B_MMP1_g NET16 N_VDD_D0_noxref_neg PFET L=6.5e-08 W=9.6e-07
+ AD=2.184e-13 AS=2.136e-13 PD=1.415e-06 PS=1.405e-06 NRD=0.236979 NRS=0.231771
+ M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=7.52e-07 SB=7.51e-07 SD=0
+ PANW1=0 PANW2=0 PANW3=1.885e-15 PANW4=3.25e-15 PANW5=3.25e-15 PANW6=6.5e-15
+ PANW7=1.3e-14 PANW8=1.3e-14 PANW9=4.121e-14 PANW10=3.9e-14
XMMP2 N_OUT_MMP2_d N_C_MMP2_g NET016 N_VDD_D0_noxref_neg PFET L=6.5e-08
+ W=9.6e-07 AD=2.2176e-13 AS=2.184e-13 PD=2.382e-06 PS=1.415e-06 NRD=0.114583
+ NRS=0.236979 M=1 NF=1 CNR_SWITCH=0 PCCRIT=0 PAR=1 PTWELL=1 SA=1.272e-06
+ SB=2.31e-07 SD=0 PANW1=0 PANW2=0 PANW3=1.885e-15 PANW4=3.25e-15 PANW5=3.25e-15
+ PANW6=6.5e-15 PANW7=1.3e-14 PANW8=1.3e-14 PANW9=4.121e-14 PANW10=1.014e-13
c_167 NET16 0 1.35129e-19
c_170 NET016 0 1.35129e-19
*
.include "/home/012/k/kt/ktd170030/cad/gf65/NOR3_PEX/nor3.pex.sp.NOR3.pxi"
*
.ends
*
*
